// rom.v
// to be included from the top module at the comple

`define MEM(x, y) {mem_hi[(x)/2], mem_lo[(x)/2]}=y

initial
begin
`MEM('o001000, 16'o012706);
`MEM('o001002, 16'o010000);
`MEM('o001004, 16'o004767);
`MEM('o001006, 16'o000122);
`MEM('o001010, 16'o010546);
`MEM('o001012, 16'o010605);
`MEM('o001014, 16'o000240);
`MEM('o001016, 16'o016700);
`MEM('o001020, 16'o000156);
`MEM('o001022, 16'o011000);
`MEM('o001024, 16'o042700);
`MEM('o001026, 16'o177577);
`MEM('o001030, 16'o005700);
`MEM('o001032, 16'o001771);
`MEM('o001034, 16'o016700);
`MEM('o001036, 16'o000140);
`MEM('o001040, 16'o016560);
`MEM('o001042, 16'o000004);
`MEM('o001044, 16'o000002);
`MEM('o001046, 16'o000240);
`MEM('o001050, 16'o012605);
`MEM('o001052, 16'o000207);
`MEM('o001054, 16'o010546);
`MEM('o001056, 16'o010605);
`MEM('o001060, 16'o000415);
`MEM('o001062, 16'o016500);
`MEM('o001064, 16'o000004);
`MEM('o001066, 16'o010001);
`MEM('o001070, 16'o005201);
`MEM('o001072, 16'o010165);
`MEM('o001074, 16'o000004);
`MEM('o001076, 16'o111000);
`MEM('o001100, 16'o110000);
`MEM('o001102, 16'o010046);
`MEM('o001104, 16'o004767);
`MEM('o001106, 16'o177700);
`MEM('o001110, 16'o062706);
`MEM('o001112, 16'o000002);
`MEM('o001114, 16'o117500);
`MEM('o001116, 16'o000004);
`MEM('o001120, 16'o105700);
`MEM('o001122, 16'o001357);
`MEM('o001124, 16'o005000);
`MEM('o001126, 16'o012605);
`MEM('o001130, 16'o000207);
`MEM('o001132, 16'o010546);
`MEM('o001134, 16'o010605);
`MEM('o001136, 16'o012746);
`MEM('o001140, 16'o001202);
`MEM('o001142, 16'o004767);
`MEM('o001144, 16'o177706);
`MEM('o001146, 16'o062706);
`MEM('o001150, 16'o000002);
`MEM('o001152, 16'o000777);
`MEM('o001154, 16'o000000);
`MEM('o001156, 16'o000000);
`MEM('o001160, 16'o000000);
`MEM('o001162, 16'o000000);
`MEM('o001164, 16'o000000);
`MEM('o001166, 16'o000000);
`MEM('o001170, 16'o000000);
`MEM('o001172, 16'o000000);
`MEM('o001174, 16'o000000);
`MEM('o001176, 16'o000000);
`MEM('o001200, 16'o177564);
`MEM('o001202, 16'o062510);
`MEM('o001204, 16'o066154);
`MEM('o001206, 16'o026157);
`MEM('o001210, 16'o053440);
`MEM('o001212, 16'o071157);
`MEM('o001214, 16'o062154);
`MEM('o001216, 16'o005041);
`MEM('o001220, 16'o000015);
`MEM('o001222, 16'o000000);
`MEM('o001224, 16'o000000);
`MEM('o001226, 16'o000000);
`MEM('o001230, 16'o000000);
`MEM('o001232, 16'o000000);
`MEM('o001234, 16'o000000);
`MEM('o001236, 16'o000000);
`MEM('o001240, 16'o000000);
`MEM('o001242, 16'o000000);
`MEM('o001244, 16'o000000);
`MEM('o001246, 16'o000000);
`MEM('o001250, 16'o000000);
`MEM('o001252, 16'o000000);
`MEM('o001254, 16'o000000);
`MEM('o001256, 16'o000000);
`MEM('o001260, 16'o000000);
`MEM('o001262, 16'o000000);
`MEM('o001264, 16'o000000);
`MEM('o001266, 16'o000000);
`MEM('o001270, 16'o000000);
`MEM('o001272, 16'o000000);
`MEM('o001274, 16'o000000);
`MEM('o001276, 16'o000000);
`MEM('o001300, 16'o000000);
`MEM('o001302, 16'o000004);
`MEM('o001304, 16'o000002);
`MEM('o001306, 16'o001000);
`MEM('o001310, 16'o000000);
`MEM('o001312, 16'o000014);
`MEM('o001314, 16'o000042);
`MEM('o001316, 16'o001000);
`MEM('o001320, 16'o000000);
`MEM('o001322, 16'o000022);
`MEM('o001324, 16'o000042);
`MEM('o001326, 16'o001132);
`MEM('o001330, 16'o000000);
`MEM('o001332, 16'o000032);
`MEM('o001334, 16'o000002);
`MEM('o001336, 16'o001010);
`MEM('o001340, 16'o000000);
`MEM('o001342, 16'o000042);
`MEM('o001344, 16'o000003);
`MEM('o001346, 16'o001200);
`MEM('o001350, 16'o000000);
`MEM('o001352, 16'o000051);
`MEM('o001354, 16'o000042);
`MEM('o001356, 16'o001010);
`MEM('o001360, 16'o000000);
`MEM('o001362, 16'o000062);
`MEM('o001364, 16'o000042);
`MEM('o001366, 16'o001054);
`MEM('o001370, 16'o000000);
`MEM('o001372, 16'o000070);
`MEM('o001374, 16'o072163);
`MEM('o001376, 16'o071141);
`MEM('o001400, 16'o027164);
`MEM('o001402, 16'o000157);
`MEM('o001404, 16'o072163);
`MEM('o001406, 16'o071141);
`MEM('o001410, 16'o000164);
`MEM('o001412, 16'o061537);
`MEM('o001414, 16'o072163);
`MEM('o001416, 16'o071141);
`MEM('o001420, 16'o000164);
`MEM('o001422, 16'o062550);
`MEM('o001424, 16'o066154);
`MEM('o001426, 16'o027157);
`MEM('o001430, 16'o000157);
`MEM('o001432, 16'o070137);
`MEM('o001434, 16'o066153);
`MEM('o001436, 16'o030461);
`MEM('o001440, 16'o057400);
`MEM('o001442, 16'o072560);
`MEM('o001444, 16'o061564);
`MEM('o001446, 16'o060550);
`MEM('o001450, 16'o000162);
`MEM('o001452, 16'o070137);
`MEM('o001454, 16'o072165);
`MEM('o001456, 16'o000163);
`MEM('o001460, 16'o000000);
`MEM('o001462, 16'o000000);
`MEM('o001464, 16'o000000);
`MEM('o001466, 16'o000000);
`MEM('o001470, 16'o000000);
`MEM('o001472, 16'o000000);
`MEM('o001474, 16'o000000);
`MEM('o001476, 16'o000000);
`MEM('o001500, 16'o000000);
`MEM('o001502, 16'o000000);
`MEM('o001504, 16'o000000);
`MEM('o001506, 16'o000000);
`MEM('o001510, 16'o000000);
`MEM('o001512, 16'o000000);
`MEM('o001514, 16'o000000);
`MEM('o001516, 16'o000000);
`MEM('o001520, 16'o000000);
`MEM('o001522, 16'o000000);
`MEM('o001524, 16'o000000);
`MEM('o001526, 16'o000000);
`MEM('o001530, 16'o000000);
`MEM('o001532, 16'o000000);
`MEM('o001534, 16'o000000);
`MEM('o001536, 16'o000000);
`MEM('o001540, 16'o000000);
`MEM('o001542, 16'o000000);
`MEM('o001544, 16'o000000);
`MEM('o001546, 16'o000000);
`MEM('o001550, 16'o000000);
`MEM('o001552, 16'o000000);
`MEM('o001554, 16'o000000);
`MEM('o001556, 16'o000000);
`MEM('o001560, 16'o000000);
`MEM('o001562, 16'o000000);
`MEM('o001564, 16'o000000);
`MEM('o001566, 16'o000000);
`MEM('o001570, 16'o000000);
`MEM('o001572, 16'o000000);
`MEM('o001574, 16'o000000);
`MEM('o001576, 16'o000000);
`MEM('o001600, 16'o000000);
`MEM('o001602, 16'o000000);
`MEM('o001604, 16'o000000);
`MEM('o001606, 16'o000000);
`MEM('o001610, 16'o000000);
`MEM('o001612, 16'o000000);
`MEM('o001614, 16'o000000);
`MEM('o001616, 16'o000000);
`MEM('o001620, 16'o000000);
`MEM('o001622, 16'o000000);
`MEM('o001624, 16'o000000);
`MEM('o001626, 16'o000000);
`MEM('o001630, 16'o000000);
`MEM('o001632, 16'o000000);
`MEM('o001634, 16'o000000);
`MEM('o001636, 16'o000000);
`MEM('o001640, 16'o000000);
`MEM('o001642, 16'o000000);
`MEM('o001644, 16'o000000);
`MEM('o001646, 16'o000000);
`MEM('o001650, 16'o000000);
`MEM('o001652, 16'o000000);
`MEM('o001654, 16'o000000);
`MEM('o001656, 16'o000000);
`MEM('o001660, 16'o000000);
`MEM('o001662, 16'o000000);
`MEM('o001664, 16'o000000);
`MEM('o001666, 16'o000000);
`MEM('o001670, 16'o000000);
`MEM('o001672, 16'o000000);
`MEM('o001674, 16'o000000);
`MEM('o001676, 16'o000000);
`MEM('o001700, 16'o000000);
`MEM('o001702, 16'o000000);
`MEM('o001704, 16'o000000);
`MEM('o001706, 16'o000000);
`MEM('o001710, 16'o000000);
`MEM('o001712, 16'o000000);
`MEM('o001714, 16'o000000);
`MEM('o001716, 16'o000000);
`MEM('o001720, 16'o000000);
`MEM('o001722, 16'o000000);
`MEM('o001724, 16'o000000);
`MEM('o001726, 16'o000000);
`MEM('o001730, 16'o000000);
`MEM('o001732, 16'o000000);
`MEM('o001734, 16'o000000);
`MEM('o001736, 16'o000000);
`MEM('o001740, 16'o000000);
`MEM('o001742, 16'o000000);
`MEM('o001744, 16'o000000);
`MEM('o001746, 16'o000000);
`MEM('o001750, 16'o000000);
`MEM('o001752, 16'o000000);
`MEM('o001754, 16'o000000);
`MEM('o001756, 16'o000000);
`MEM('o001760, 16'o000000);
`MEM('o001762, 16'o000000);
`MEM('o001764, 16'o000000);
`MEM('o001766, 16'o000000);
`MEM('o001770, 16'o000000);
`MEM('o001772, 16'o000000);
`MEM('o001774, 16'o000000);
`MEM('o001776, 16'o000000);
end
