// rom.v
// to be included from the top module at the comple

`define MEM(x, y) {mem_hi[(x)/2], mem_lo[(x)/2]}=y

initial
begin
`MEM('o001000, 16'o012706);
`MEM('o001002, 16'o001000);
`MEM('o001004, 16'o004767);
`MEM('o001006, 16'o017020);
`MEM('o001010, 16'o010546);
`MEM('o001012, 16'o010605);
`MEM('o001014, 16'o000240);
`MEM('o001016, 16'o012700);
`MEM('o001020, 16'o177564);
`MEM('o001022, 16'o111000);
`MEM('o001024, 16'o105700);
`MEM('o001026, 16'o002373);
`MEM('o001030, 16'o012700);
`MEM('o001032, 16'o177566);
`MEM('o001034, 16'o016501);
`MEM('o001036, 16'o000004);
`MEM('o001040, 16'o110110);
`MEM('o001042, 16'o000240);
`MEM('o001044, 16'o012605);
`MEM('o001046, 16'o000207);
`MEM('o001050, 16'o010546);
`MEM('o001052, 16'o010605);
`MEM('o001054, 16'o000240);
`MEM('o001056, 16'o012700);
`MEM('o001060, 16'o177560);
`MEM('o001062, 16'o111000);
`MEM('o001064, 16'o105700);
`MEM('o001066, 16'o002373);
`MEM('o001070, 16'o012700);
`MEM('o001072, 16'o177562);
`MEM('o001074, 16'o111000);
`MEM('o001076, 16'o042700);
`MEM('o001100, 16'o177400);
`MEM('o001102, 16'o012605);
`MEM('o001104, 16'o000207);
`MEM('o001106, 16'o010546);
`MEM('o001110, 16'o010605);
`MEM('o001112, 16'o012700);
`MEM('o001114, 16'o177560);
`MEM('o001116, 16'o111000);
`MEM('o001120, 16'o042700);
`MEM('o001122, 16'o177400);
`MEM('o001124, 16'o072027);
`MEM('o001126, 16'o000007);
`MEM('o001130, 16'o042700);
`MEM('o001132, 16'o177400);
`MEM('o001134, 16'o012605);
`MEM('o001136, 16'o000207);
`MEM('o001140, 16'o010546);
`MEM('o001142, 16'o010605);
`MEM('o001144, 16'o012746);
`MEM('o001146, 16'o000015);
`MEM('o001150, 16'o004767);
`MEM('o001152, 16'o177634);
`MEM('o001154, 16'o062706);
`MEM('o001156, 16'o000002);
`MEM('o001160, 16'o012746);
`MEM('o001162, 16'o000012);
`MEM('o001164, 16'o004767);
`MEM('o001166, 16'o177620);
`MEM('o001170, 16'o062706);
`MEM('o001172, 16'o000002);
`MEM('o001174, 16'o000240);
`MEM('o001176, 16'o012605);
`MEM('o001200, 16'o000207);
`MEM('o001202, 16'o010546);
`MEM('o001204, 16'o010605);
`MEM('o001206, 16'o000414);
`MEM('o001210, 16'o005000);
`MEM('o001212, 16'o156500);
`MEM('o001214, 16'o000010);
`MEM('o001216, 16'o066500);
`MEM('o001220, 16'o000006);
`MEM('o001222, 16'o111000);
`MEM('o001224, 16'o126500);
`MEM('o001226, 16'o000004);
`MEM('o001230, 16'o001003);
`MEM('o001232, 16'o112700);
`MEM('o001234, 16'o000001);
`MEM('o001236, 16'o000411);
`MEM('o001240, 16'o116500);
`MEM('o001242, 16'o000010);
`MEM('o001244, 16'o110001);
`MEM('o001246, 16'o105301);
`MEM('o001250, 16'o110165);
`MEM('o001252, 16'o000010);
`MEM('o001254, 16'o105700);
`MEM('o001256, 16'o001354);
`MEM('o001260, 16'o105000);
`MEM('o001262, 16'o012605);
`MEM('o001264, 16'o000207);
`MEM('o001266, 16'o010546);
`MEM('o001270, 16'o010605);
`MEM('o001272, 16'o126527);
`MEM('o001274, 16'o000004);
`MEM('o001276, 16'o000172);
`MEM('o001300, 16'o003011);
`MEM('o001302, 16'o126527);
`MEM('o001304, 16'o000004);
`MEM('o001306, 16'o000140);
`MEM('o001310, 16'o003405);
`MEM('o001312, 16'o116500);
`MEM('o001314, 16'o000004);
`MEM('o001316, 16'o062700);
`MEM('o001320, 16'o177740);
`MEM('o001322, 16'o000402);
`MEM('o001324, 16'o116500);
`MEM('o001326, 16'o000004);
`MEM('o001330, 16'o012605);
`MEM('o001332, 16'o000207);
`MEM('o001334, 16'o010546);
`MEM('o001336, 16'o010605);
`MEM('o001340, 16'o126527);
`MEM('o001342, 16'o000004);
`MEM('o001344, 16'o000037);
`MEM('o001346, 16'o003407);
`MEM('o001350, 16'o126527);
`MEM('o001352, 16'o000004);
`MEM('o001354, 16'o000177);
`MEM('o001356, 16'o001403);
`MEM('o001360, 16'o012700);
`MEM('o001362, 16'o000001);
`MEM('o001364, 16'o000401);
`MEM('o001366, 16'o005000);
`MEM('o001370, 16'o012605);
`MEM('o001372, 16'o000207);
`MEM('o001374, 16'o010546);
`MEM('o001376, 16'o010605);
`MEM('o001400, 16'o126527);
`MEM('o001402, 16'o000004);
`MEM('o001404, 16'o000040);
`MEM('o001406, 16'o001410);
`MEM('o001410, 16'o126527);
`MEM('o001412, 16'o000004);
`MEM('o001414, 16'o000015);
`MEM('o001416, 16'o003007);
`MEM('o001420, 16'o126527);
`MEM('o001422, 16'o000004);
`MEM('o001424, 16'o000010);
`MEM('o001426, 16'o003403);
`MEM('o001430, 16'o012700);
`MEM('o001432, 16'o000001);
`MEM('o001434, 16'o000401);
`MEM('o001436, 16'o005000);
`MEM('o001440, 16'o012605);
`MEM('o001442, 16'o000207);
`MEM('o001444, 16'o010546);
`MEM('o001446, 16'o010605);
`MEM('o001450, 16'o126527);
`MEM('o001452, 16'o000004);
`MEM('o001454, 16'o000071);
`MEM('o001456, 16'o003007);
`MEM('o001460, 16'o126527);
`MEM('o001462, 16'o000004);
`MEM('o001464, 16'o000057);
`MEM('o001466, 16'o003403);
`MEM('o001470, 16'o012700);
`MEM('o001472, 16'o000001);
`MEM('o001474, 16'o000401);
`MEM('o001476, 16'o005000);
`MEM('o001500, 16'o012605);
`MEM('o001502, 16'o000207);
`MEM('o001504, 16'o010546);
`MEM('o001506, 16'o010605);
`MEM('o001510, 16'o126527);
`MEM('o001512, 16'o000004);
`MEM('o001514, 16'o000172);
`MEM('o001516, 16'o003004);
`MEM('o001520, 16'o126527);
`MEM('o001522, 16'o000004);
`MEM('o001524, 16'o000140);
`MEM('o001526, 16'o003010);
`MEM('o001530, 16'o126527);
`MEM('o001532, 16'o000004);
`MEM('o001534, 16'o000132);
`MEM('o001536, 16'o003007);
`MEM('o001540, 16'o126527);
`MEM('o001542, 16'o000004);
`MEM('o001544, 16'o000100);
`MEM('o001546, 16'o003403);
`MEM('o001550, 16'o012700);
`MEM('o001552, 16'o000001);
`MEM('o001554, 16'o000401);
`MEM('o001556, 16'o005000);
`MEM('o001560, 16'o012605);
`MEM('o001562, 16'o000207);
`MEM('o001564, 16'o010546);
`MEM('o001566, 16'o010605);
`MEM('o001570, 16'o000415);
`MEM('o001572, 16'o016500);
`MEM('o001574, 16'o000004);
`MEM('o001576, 16'o010001);
`MEM('o001600, 16'o005201);
`MEM('o001602, 16'o010165);
`MEM('o001604, 16'o000004);
`MEM('o001606, 16'o111000);
`MEM('o001610, 16'o110000);
`MEM('o001612, 16'o010046);
`MEM('o001614, 16'o004767);
`MEM('o001616, 16'o177170);
`MEM('o001620, 16'o062706);
`MEM('o001622, 16'o000002);
`MEM('o001624, 16'o117500);
`MEM('o001626, 16'o000004);
`MEM('o001630, 16'o105700);
`MEM('o001632, 16'o001357);
`MEM('o001634, 16'o000240);
`MEM('o001636, 16'o000240);
`MEM('o001640, 16'o012605);
`MEM('o001642, 16'o000207);
`MEM('o001644, 16'o010546);
`MEM('o001646, 16'o010605);
`MEM('o001650, 16'o062706);
`MEM('o001652, 16'o177776);
`MEM('o001654, 16'o105065);
`MEM('o001656, 16'o177776);
`MEM('o001660, 16'o000511);
`MEM('o001662, 16'o126527);
`MEM('o001664, 16'o177777);
`MEM('o001666, 16'o000011);
`MEM('o001670, 16'o001003);
`MEM('o001672, 16'o112765);
`MEM('o001674, 16'o000040);
`MEM('o001676, 16'o177777);
`MEM('o001700, 16'o126527);
`MEM('o001702, 16'o177777);
`MEM('o001704, 16'o000010);
`MEM('o001706, 16'o001404);
`MEM('o001710, 16'o126527);
`MEM('o001712, 16'o177777);
`MEM('o001714, 16'o000177);
`MEM('o001716, 16'o001034);
`MEM('o001720, 16'o105765);
`MEM('o001722, 16'o177776);
`MEM('o001724, 16'o001431);
`MEM('o001726, 16'o116500);
`MEM('o001730, 16'o177776);
`MEM('o001732, 16'o110001);
`MEM('o001734, 16'o105301);
`MEM('o001736, 16'o110165);
`MEM('o001740, 16'o177776);
`MEM('o001742, 16'o012746);
`MEM('o001744, 16'o000010);
`MEM('o001746, 16'o004767);
`MEM('o001750, 16'o177036);
`MEM('o001752, 16'o062706);
`MEM('o001754, 16'o000002);
`MEM('o001756, 16'o012746);
`MEM('o001760, 16'o000040);
`MEM('o001762, 16'o004767);
`MEM('o001764, 16'o177022);
`MEM('o001766, 16'o062706);
`MEM('o001770, 16'o000002);
`MEM('o001772, 16'o012746);
`MEM('o001774, 16'o000010);
`MEM('o001776, 16'o004767);
`MEM('o002000, 16'o177006);
`MEM('o002002, 16'o062706);
`MEM('o002004, 16'o000002);
`MEM('o002006, 16'o000436);
`MEM('o002010, 16'o116546);
`MEM('o002012, 16'o177777);
`MEM('o002014, 16'o004767);
`MEM('o002016, 16'o177314);
`MEM('o002020, 16'o062706);
`MEM('o002022, 16'o000002);
`MEM('o002024, 16'o105700);
`MEM('o002026, 16'o001426);
`MEM('o002030, 16'o126527);
`MEM('o002032, 16'o177776);
`MEM('o002034, 16'o000116);
`MEM('o002036, 16'o101022);
`MEM('o002040, 16'o116500);
`MEM('o002042, 16'o177776);
`MEM('o002044, 16'o110001);
`MEM('o002046, 16'o105201);
`MEM('o002050, 16'o110165);
`MEM('o002052, 16'o177776);
`MEM('o002054, 16'o042700);
`MEM('o002056, 16'o177400);
`MEM('o002060, 16'o116560);
`MEM('o002062, 16'o177777);
`MEM('o002064, 16'o021540);
`MEM('o002066, 16'o116500);
`MEM('o002070, 16'o177777);
`MEM('o002072, 16'o010046);
`MEM('o002074, 16'o004767);
`MEM('o002076, 16'o176710);
`MEM('o002100, 16'o062706);
`MEM('o002102, 16'o000002);
`MEM('o002104, 16'o004767);
`MEM('o002106, 16'o176740);
`MEM('o002110, 16'o110065);
`MEM('o002112, 16'o177777);
`MEM('o002114, 16'o126527);
`MEM('o002116, 16'o177777);
`MEM('o002120, 16'o000015);
`MEM('o002122, 16'o001257);
`MEM('o002124, 16'o004767);
`MEM('o002126, 16'o177010);
`MEM('o002130, 16'o005000);
`MEM('o002132, 16'o156500);
`MEM('o002134, 16'o177776);
`MEM('o002136, 16'o105060);
`MEM('o002140, 16'o021540);
`MEM('o002142, 16'o105765);
`MEM('o002144, 16'o177776);
`MEM('o002146, 16'o001426);
`MEM('o002150, 16'o000240);
`MEM('o002152, 16'o105365);
`MEM('o002154, 16'o177776);
`MEM('o002156, 16'o005000);
`MEM('o002160, 16'o156500);
`MEM('o002162, 16'o177776);
`MEM('o002164, 16'o116000);
`MEM('o002166, 16'o021540);
`MEM('o002170, 16'o110046);
`MEM('o002172, 16'o004767);
`MEM('o002174, 16'o177176);
`MEM('o002176, 16'o062706);
`MEM('o002200, 16'o000002);
`MEM('o002202, 16'o105700);
`MEM('o002204, 16'o001362);
`MEM('o002206, 16'o105265);
`MEM('o002210, 16'o177776);
`MEM('o002212, 16'o005000);
`MEM('o002214, 16'o156500);
`MEM('o002216, 16'o177776);
`MEM('o002220, 16'o105060);
`MEM('o002222, 16'o021540);
`MEM('o002224, 16'o000240);
`MEM('o002226, 16'o010506);
`MEM('o002230, 16'o012605);
`MEM('o002232, 16'o000207);
`MEM('o002234, 16'o010546);
`MEM('o002236, 16'o010605);
`MEM('o002240, 16'o062706);
`MEM('o002242, 16'o177776);
`MEM('o002244, 16'o005765);
`MEM('o002246, 16'o000004);
`MEM('o002250, 16'o002006);
`MEM('o002252, 16'o112765);
`MEM('o002254, 16'o000001);
`MEM('o002256, 16'o177776);
`MEM('o002260, 16'o005465);
`MEM('o002262, 16'o000004);
`MEM('o002264, 16'o000402);
`MEM('o002266, 16'o105065);
`MEM('o002270, 16'o177776);
`MEM('o002272, 16'o105067);
`MEM('o002274, 16'o017250);
`MEM('o002276, 16'o112765);
`MEM('o002300, 16'o000006);
`MEM('o002302, 16'o177777);
`MEM('o002304, 16'o016500);
`MEM('o002306, 16'o000004);
`MEM('o002310, 16'o010001);
`MEM('o002312, 16'o006700);
`MEM('o002314, 16'o071027);
`MEM('o002316, 16'o000012);
`MEM('o002320, 16'o010100);
`MEM('o002322, 16'o062700);
`MEM('o002324, 16'o000060);
`MEM('o002326, 16'o110001);
`MEM('o002330, 16'o105365);
`MEM('o002332, 16'o177777);
`MEM('o002334, 16'o005000);
`MEM('o002336, 16'o156500);
`MEM('o002340, 16'o177777);
`MEM('o002342, 16'o110160);
`MEM('o002344, 16'o021540);
`MEM('o002346, 16'o016500);
`MEM('o002350, 16'o000004);
`MEM('o002352, 16'o010001);
`MEM('o002354, 16'o006700);
`MEM('o002356, 16'o071027);
`MEM('o002360, 16'o000012);
`MEM('o002362, 16'o010065);
`MEM('o002364, 16'o000004);
`MEM('o002366, 16'o005765);
`MEM('o002370, 16'o000004);
`MEM('o002372, 16'o003344);
`MEM('o002374, 16'o105765);
`MEM('o002376, 16'o177776);
`MEM('o002400, 16'o001424);
`MEM('o002402, 16'o105365);
`MEM('o002404, 16'o177777);
`MEM('o002406, 16'o005000);
`MEM('o002410, 16'o156500);
`MEM('o002412, 16'o177777);
`MEM('o002414, 16'o112760);
`MEM('o002416, 16'o000055);
`MEM('o002420, 16'o021540);
`MEM('o002422, 16'o000413);
`MEM('o002424, 16'o012746);
`MEM('o002426, 16'o000040);
`MEM('o002430, 16'o004767);
`MEM('o002432, 16'o176354);
`MEM('o002434, 16'o062706);
`MEM('o002436, 16'o000002);
`MEM('o002440, 16'o016500);
`MEM('o002442, 16'o000006);
`MEM('o002444, 16'o005300);
`MEM('o002446, 16'o010065);
`MEM('o002450, 16'o000006);
`MEM('o002452, 16'o005000);
`MEM('o002454, 16'o156500);
`MEM('o002456, 16'o177777);
`MEM('o002460, 16'o012701);
`MEM('o002462, 16'o000006);
`MEM('o002464, 16'o160001);
`MEM('o002466, 16'o026501);
`MEM('o002470, 16'o000006);
`MEM('o002472, 16'o003354);
`MEM('o002474, 16'o005000);
`MEM('o002476, 16'o156500);
`MEM('o002500, 16'o177777);
`MEM('o002502, 16'o062700);
`MEM('o002504, 16'o021540);
`MEM('o002506, 16'o010046);
`MEM('o002510, 16'o004767);
`MEM('o002512, 16'o177050);
`MEM('o002514, 16'o062706);
`MEM('o002516, 16'o000002);
`MEM('o002520, 16'o000240);
`MEM('o002522, 16'o010506);
`MEM('o002524, 16'o012605);
`MEM('o002526, 16'o000207);
`MEM('o002530, 16'o010246);
`MEM('o002532, 16'o010546);
`MEM('o002534, 16'o010605);
`MEM('o002536, 16'o062706);
`MEM('o002540, 16'o177770);
`MEM('o002542, 16'o105065);
`MEM('o002544, 16'o177775);
`MEM('o002546, 16'o000515);
`MEM('o002550, 16'o126527);
`MEM('o002552, 16'o177773);
`MEM('o002554, 16'o000010);
`MEM('o002556, 16'o001404);
`MEM('o002560, 16'o126527);
`MEM('o002562, 16'o177773);
`MEM('o002564, 16'o000177);
`MEM('o002566, 16'o001034);
`MEM('o002570, 16'o105765);
`MEM('o002572, 16'o177775);
`MEM('o002574, 16'o001431);
`MEM('o002576, 16'o116500);
`MEM('o002600, 16'o177775);
`MEM('o002602, 16'o110001);
`MEM('o002604, 16'o105301);
`MEM('o002606, 16'o110165);
`MEM('o002610, 16'o177775);
`MEM('o002612, 16'o012746);
`MEM('o002614, 16'o000010);
`MEM('o002616, 16'o004767);
`MEM('o002620, 16'o176166);
`MEM('o002622, 16'o062706);
`MEM('o002624, 16'o000002);
`MEM('o002626, 16'o012746);
`MEM('o002630, 16'o000040);
`MEM('o002632, 16'o004767);
`MEM('o002634, 16'o176152);
`MEM('o002636, 16'o062706);
`MEM('o002640, 16'o000002);
`MEM('o002642, 16'o012746);
`MEM('o002644, 16'o000010);
`MEM('o002646, 16'o004767);
`MEM('o002650, 16'o176136);
`MEM('o002652, 16'o062706);
`MEM('o002654, 16'o000002);
`MEM('o002656, 16'o000451);
`MEM('o002660, 16'o105765);
`MEM('o002662, 16'o177775);
`MEM('o002664, 16'o001010);
`MEM('o002666, 16'o126527);
`MEM('o002670, 16'o177773);
`MEM('o002672, 16'o000053);
`MEM('o002674, 16'o001420);
`MEM('o002676, 16'o126527);
`MEM('o002700, 16'o177773);
`MEM('o002702, 16'o000055);
`MEM('o002704, 16'o001414);
`MEM('o002706, 16'o126527);
`MEM('o002710, 16'o177775);
`MEM('o002712, 16'o000005);
`MEM('o002714, 16'o101032);
`MEM('o002716, 16'o116546);
`MEM('o002720, 16'o177773);
`MEM('o002722, 16'o004767);
`MEM('o002724, 16'o176516);
`MEM('o002726, 16'o062706);
`MEM('o002730, 16'o000002);
`MEM('o002732, 16'o105700);
`MEM('o002734, 16'o001422);
`MEM('o002736, 16'o116500);
`MEM('o002740, 16'o177775);
`MEM('o002742, 16'o110002);
`MEM('o002744, 16'o105202);
`MEM('o002746, 16'o110265);
`MEM('o002750, 16'o177775);
`MEM('o002752, 16'o042700);
`MEM('o002754, 16'o177400);
`MEM('o002756, 16'o116560);
`MEM('o002760, 16'o177773);
`MEM('o002762, 16'o021540);
`MEM('o002764, 16'o116500);
`MEM('o002766, 16'o177773);
`MEM('o002770, 16'o010046);
`MEM('o002772, 16'o004767);
`MEM('o002774, 16'o176012);
`MEM('o002776, 16'o062706);
`MEM('o003000, 16'o000002);
`MEM('o003002, 16'o004767);
`MEM('o003004, 16'o176042);
`MEM('o003006, 16'o110065);
`MEM('o003010, 16'o177773);
`MEM('o003012, 16'o126527);
`MEM('o003014, 16'o177773);
`MEM('o003016, 16'o000015);
`MEM('o003020, 16'o001253);
`MEM('o003022, 16'o004767);
`MEM('o003024, 16'o176112);
`MEM('o003026, 16'o005000);
`MEM('o003030, 16'o156500);
`MEM('o003032, 16'o177775);
`MEM('o003034, 16'o105060);
`MEM('o003036, 16'o021540);
`MEM('o003040, 16'o116700);
`MEM('o003042, 16'o016474);
`MEM('o003044, 16'o110000);
`MEM('o003046, 16'o020027);
`MEM('o003050, 16'o000053);
`MEM('o003052, 16'o001412);
`MEM('o003054, 16'o020027);
`MEM('o003056, 16'o000055);
`MEM('o003060, 16'o001015);
`MEM('o003062, 16'o112765);
`MEM('o003064, 16'o000001);
`MEM('o003066, 16'o177774);
`MEM('o003070, 16'o112765);
`MEM('o003072, 16'o000001);
`MEM('o003074, 16'o177775);
`MEM('o003076, 16'o000413);
`MEM('o003100, 16'o105065);
`MEM('o003102, 16'o177774);
`MEM('o003104, 16'o112765);
`MEM('o003106, 16'o000001);
`MEM('o003110, 16'o177775);
`MEM('o003112, 16'o000405);
`MEM('o003114, 16'o105065);
`MEM('o003116, 16'o177774);
`MEM('o003120, 16'o105065);
`MEM('o003122, 16'o177775);
`MEM('o003124, 16'o000240);
`MEM('o003126, 16'o005065);
`MEM('o003130, 16'o177776);
`MEM('o003132, 16'o005065);
`MEM('o003134, 16'o177770);
`MEM('o003136, 16'o000443);
`MEM('o003140, 16'o016501);
`MEM('o003142, 16'o177776);
`MEM('o003144, 16'o010100);
`MEM('o003146, 16'o006300);
`MEM('o003150, 16'o006300);
`MEM('o003152, 16'o060100);
`MEM('o003154, 16'o006300);
`MEM('o003156, 16'o010001);
`MEM('o003160, 16'o116500);
`MEM('o003162, 16'o177775);
`MEM('o003164, 16'o110002);
`MEM('o003166, 16'o105202);
`MEM('o003170, 16'o110265);
`MEM('o003172, 16'o177775);
`MEM('o003174, 16'o042700);
`MEM('o003176, 16'o177400);
`MEM('o003200, 16'o116000);
`MEM('o003202, 16'o021540);
`MEM('o003204, 16'o110000);
`MEM('o003206, 16'o060100);
`MEM('o003210, 16'o012701);
`MEM('o003212, 16'o177720);
`MEM('o003214, 16'o060001);
`MEM('o003216, 16'o010165);
`MEM('o003220, 16'o177770);
`MEM('o003222, 16'o026565);
`MEM('o003224, 16'o177776);
`MEM('o003226, 16'o177770);
`MEM('o003230, 16'o003403);
`MEM('o003232, 16'o112767);
`MEM('o003234, 16'o000002);
`MEM('o003236, 16'o015410);
`MEM('o003240, 16'o016565);
`MEM('o003242, 16'o177770);
`MEM('o003244, 16'o177776);
`MEM('o003246, 16'o005000);
`MEM('o003250, 16'o156500);
`MEM('o003252, 16'o177775);
`MEM('o003254, 16'o116000);
`MEM('o003256, 16'o021540);
`MEM('o003260, 16'o105700);
`MEM('o003262, 16'o001326);
`MEM('o003264, 16'o105765);
`MEM('o003266, 16'o177774);
`MEM('o003270, 16'o001404);
`MEM('o003272, 16'o016500);
`MEM('o003274, 16'o177776);
`MEM('o003276, 16'o005400);
`MEM('o003300, 16'o000402);
`MEM('o003302, 16'o016500);
`MEM('o003304, 16'o177776);
`MEM('o003306, 16'o010506);
`MEM('o003310, 16'o012605);
`MEM('o003312, 16'o012602);
`MEM('o003314, 16'o000207);
`MEM('o003316, 16'o010246);
`MEM('o003320, 16'o010546);
`MEM('o003322, 16'o010605);
`MEM('o003324, 16'o062706);
`MEM('o003326, 16'o177762);
`MEM('o003330, 16'o105065);
`MEM('o003332, 16'o177776);
`MEM('o003334, 16'o005065);
`MEM('o003336, 16'o177774);
`MEM('o003340, 16'o012765);
`MEM('o003342, 16'o021540);
`MEM('o003344, 16'o177770);
`MEM('o003346, 16'o000167);
`MEM('o003350, 16'o001750);
`MEM('o003352, 16'o005265);
`MEM('o003354, 16'o177770);
`MEM('o003356, 16'o117500);
`MEM('o003360, 16'o177770);
`MEM('o003362, 16'o110046);
`MEM('o003364, 16'o004767);
`MEM('o003366, 16'o176004);
`MEM('o003370, 16'o062706);
`MEM('o003372, 16'o000002);
`MEM('o003374, 16'o105700);
`MEM('o003376, 16'o001365);
`MEM('o003400, 16'o105065);
`MEM('o003402, 16'o177777);
`MEM('o003404, 16'o000502);
`MEM('o003406, 16'o005000);
`MEM('o003410, 16'o156500);
`MEM('o003412, 16'o177777);
`MEM('o003414, 16'o006300);
`MEM('o003416, 16'o062700);
`MEM('o003420, 16'o020502);
`MEM('o003422, 16'o011065);
`MEM('o003424, 16'o177774);
`MEM('o003426, 16'o016565);
`MEM('o003430, 16'o177770);
`MEM('o003432, 16'o177772);
`MEM('o003434, 16'o000404);
`MEM('o003436, 16'o005265);
`MEM('o003440, 16'o177774);
`MEM('o003442, 16'o005265);
`MEM('o003444, 16'o177772);
`MEM('o003446, 16'o117500);
`MEM('o003450, 16'o177774);
`MEM('o003452, 16'o105700);
`MEM('o003454, 16'o001413);
`MEM('o003456, 16'o117502);
`MEM('o003460, 16'o177774);
`MEM('o003462, 16'o117500);
`MEM('o003464, 16'o177772);
`MEM('o003466, 16'o110046);
`MEM('o003470, 16'o004767);
`MEM('o003472, 16'o175572);
`MEM('o003474, 16'o062706);
`MEM('o003476, 16'o000002);
`MEM('o003500, 16'o120200);
`MEM('o003502, 16'o001755);
`MEM('o003504, 16'o117500);
`MEM('o003506, 16'o177774);
`MEM('o003510, 16'o105700);
`MEM('o003512, 16'o001031);
`MEM('o003514, 16'o126527);
`MEM('o003516, 16'o177776);
`MEM('o003520, 16'o000116);
`MEM('o003522, 16'o101406);
`MEM('o003524, 16'o112767);
`MEM('o003526, 16'o000004);
`MEM('o003530, 16'o015116);
`MEM('o003532, 16'o105000);
`MEM('o003534, 16'o000167);
`MEM('o003536, 16'o001630);
`MEM('o003540, 16'o116500);
`MEM('o003542, 16'o177776);
`MEM('o003544, 16'o110001);
`MEM('o003546, 16'o105201);
`MEM('o003550, 16'o110165);
`MEM('o003552, 16'o177776);
`MEM('o003554, 16'o042700);
`MEM('o003556, 16'o177400);
`MEM('o003560, 16'o116560);
`MEM('o003562, 16'o177777);
`MEM('o003564, 16'o021660);
`MEM('o003566, 16'o016565);
`MEM('o003570, 16'o177772);
`MEM('o003572, 16'o177770);
`MEM('o003574, 16'o000412);
`MEM('o003576, 16'o116500);
`MEM('o003600, 16'o177777);
`MEM('o003602, 16'o110002);
`MEM('o003604, 16'o105202);
`MEM('o003606, 16'o110265);
`MEM('o003610, 16'o177777);
`MEM('o003612, 16'o126527);
`MEM('o003614, 16'o177777);
`MEM('o003616, 16'o000041);
`MEM('o003620, 16'o101672);
`MEM('o003622, 16'o126527);
`MEM('o003624, 16'o177777);
`MEM('o003626, 16'o000010);
`MEM('o003630, 16'o001131);
`MEM('o003632, 16'o000402);
`MEM('o003634, 16'o005265);
`MEM('o003636, 16'o177770);
`MEM('o003640, 16'o117500);
`MEM('o003642, 16'o177770);
`MEM('o003644, 16'o110046);
`MEM('o003646, 16'o004767);
`MEM('o003650, 16'o175522);
`MEM('o003652, 16'o062706);
`MEM('o003654, 16'o000002);
`MEM('o003656, 16'o105700);
`MEM('o003660, 16'o001365);
`MEM('o003662, 16'o016565);
`MEM('o003664, 16'o177770);
`MEM('o003666, 16'o177772);
`MEM('o003670, 16'o105065);
`MEM('o003672, 16'o177777);
`MEM('o003674, 16'o000406);
`MEM('o003676, 16'o116500);
`MEM('o003700, 16'o177777);
`MEM('o003702, 16'o110001);
`MEM('o003704, 16'o105201);
`MEM('o003706, 16'o110165);
`MEM('o003710, 16'o177777);
`MEM('o003712, 16'o016500);
`MEM('o003714, 16'o177772);
`MEM('o003716, 16'o010002);
`MEM('o003720, 16'o005202);
`MEM('o003722, 16'o010265);
`MEM('o003724, 16'o177772);
`MEM('o003726, 16'o111000);
`MEM('o003730, 16'o105700);
`MEM('o003732, 16'o001361);
`MEM('o003734, 16'o005000);
`MEM('o003736, 16'o156500);
`MEM('o003740, 16'o177776);
`MEM('o003742, 16'o005001);
`MEM('o003744, 16'o156501);
`MEM('o003746, 16'o177777);
`MEM('o003750, 16'o012702);
`MEM('o003752, 16'o000116);
`MEM('o003754, 16'o160102);
`MEM('o003756, 16'o020002);
`MEM('o003760, 16'o002406);
`MEM('o003762, 16'o112767);
`MEM('o003764, 16'o000004);
`MEM('o003766, 16'o014660);
`MEM('o003770, 16'o105000);
`MEM('o003772, 16'o000167);
`MEM('o003774, 16'o001372);
`MEM('o003776, 16'o116500);
`MEM('o004000, 16'o177776);
`MEM('o004002, 16'o110001);
`MEM('o004004, 16'o105201);
`MEM('o004006, 16'o110165);
`MEM('o004010, 16'o177776);
`MEM('o004012, 16'o042700);
`MEM('o004014, 16'o177400);
`MEM('o004016, 16'o116560);
`MEM('o004020, 16'o177777);
`MEM('o004022, 16'o021660);
`MEM('o004024, 16'o000421);
`MEM('o004026, 16'o016500);
`MEM('o004030, 16'o177770);
`MEM('o004032, 16'o010002);
`MEM('o004034, 16'o005202);
`MEM('o004036, 16'o010265);
`MEM('o004040, 16'o177770);
`MEM('o004042, 16'o111001);
`MEM('o004044, 16'o116500);
`MEM('o004046, 16'o177776);
`MEM('o004050, 16'o110002);
`MEM('o004052, 16'o105202);
`MEM('o004054, 16'o110265);
`MEM('o004056, 16'o177776);
`MEM('o004060, 16'o042700);
`MEM('o004062, 16'o177400);
`MEM('o004064, 16'o110160);
`MEM('o004066, 16'o021660);
`MEM('o004070, 16'o116500);
`MEM('o004072, 16'o177777);
`MEM('o004074, 16'o110001);
`MEM('o004076, 16'o105301);
`MEM('o004100, 16'o110165);
`MEM('o004102, 16'o177777);
`MEM('o004104, 16'o105700);
`MEM('o004106, 16'o001347);
`MEM('o004110, 16'o000167);
`MEM('o004112, 16'o001222);
`MEM('o004114, 16'o117500);
`MEM('o004116, 16'o177774);
`MEM('o004120, 16'o105700);
`MEM('o004122, 16'o001002);
`MEM('o004124, 16'o000167);
`MEM('o004126, 16'o001172);
`MEM('o004130, 16'o016565);
`MEM('o004132, 16'o177770);
`MEM('o004134, 16'o177772);
`MEM('o004136, 16'o117500);
`MEM('o004140, 16'o177772);
`MEM('o004142, 16'o110046);
`MEM('o004144, 16'o004767);
`MEM('o004146, 16'o175274);
`MEM('o004150, 16'o062706);
`MEM('o004152, 16'o000002);
`MEM('o004154, 16'o105700);
`MEM('o004156, 16'o001544);
`MEM('o004160, 16'o005065);
`MEM('o004162, 16'o177766);
`MEM('o004164, 16'o005065);
`MEM('o004166, 16'o177762);
`MEM('o004170, 16'o016501);
`MEM('o004172, 16'o177766);
`MEM('o004174, 16'o010100);
`MEM('o004176, 16'o006300);
`MEM('o004200, 16'o006300);
`MEM('o004202, 16'o060100);
`MEM('o004204, 16'o006300);
`MEM('o004206, 16'o010001);
`MEM('o004210, 16'o016500);
`MEM('o004212, 16'o177772);
`MEM('o004214, 16'o010002);
`MEM('o004216, 16'o005202);
`MEM('o004220, 16'o010265);
`MEM('o004222, 16'o177772);
`MEM('o004224, 16'o111000);
`MEM('o004226, 16'o110000);
`MEM('o004230, 16'o060100);
`MEM('o004232, 16'o012701);
`MEM('o004234, 16'o177720);
`MEM('o004236, 16'o060001);
`MEM('o004240, 16'o010165);
`MEM('o004242, 16'o177762);
`MEM('o004244, 16'o026565);
`MEM('o004246, 16'o177766);
`MEM('o004250, 16'o177762);
`MEM('o004252, 16'o003406);
`MEM('o004254, 16'o112767);
`MEM('o004256, 16'o000002);
`MEM('o004260, 16'o014366);
`MEM('o004262, 16'o105000);
`MEM('o004264, 16'o000167);
`MEM('o004266, 16'o001100);
`MEM('o004270, 16'o016565);
`MEM('o004272, 16'o177762);
`MEM('o004274, 16'o177766);
`MEM('o004276, 16'o117500);
`MEM('o004300, 16'o177772);
`MEM('o004302, 16'o110046);
`MEM('o004304, 16'o004767);
`MEM('o004306, 16'o175134);
`MEM('o004310, 16'o062706);
`MEM('o004312, 16'o000002);
`MEM('o004314, 16'o105700);
`MEM('o004316, 16'o001324);
`MEM('o004320, 16'o126527);
`MEM('o004322, 16'o177776);
`MEM('o004324, 16'o000114);
`MEM('o004326, 16'o101406);
`MEM('o004330, 16'o112767);
`MEM('o004332, 16'o000004);
`MEM('o004334, 16'o014312);
`MEM('o004336, 16'o105000);
`MEM('o004340, 16'o000167);
`MEM('o004342, 16'o001024);
`MEM('o004344, 16'o116500);
`MEM('o004346, 16'o177776);
`MEM('o004350, 16'o110002);
`MEM('o004352, 16'o105202);
`MEM('o004354, 16'o110265);
`MEM('o004356, 16'o177776);
`MEM('o004360, 16'o042700);
`MEM('o004362, 16'o177400);
`MEM('o004364, 16'o112760);
`MEM('o004366, 16'o000042);
`MEM('o004370, 16'o021660);
`MEM('o004372, 16'o116500);
`MEM('o004374, 16'o177776);
`MEM('o004376, 16'o110001);
`MEM('o004400, 16'o105201);
`MEM('o004402, 16'o110165);
`MEM('o004404, 16'o177776);
`MEM('o004406, 16'o042700);
`MEM('o004410, 16'o177400);
`MEM('o004412, 16'o016501);
`MEM('o004414, 16'o177766);
`MEM('o004416, 16'o110160);
`MEM('o004420, 16'o021660);
`MEM('o004422, 16'o016501);
`MEM('o004424, 16'o177766);
`MEM('o004426, 16'o072127);
`MEM('o004430, 16'o177770);
`MEM('o004432, 16'o116500);
`MEM('o004434, 16'o177776);
`MEM('o004436, 16'o110002);
`MEM('o004440, 16'o105202);
`MEM('o004442, 16'o110265);
`MEM('o004444, 16'o177776);
`MEM('o004446, 16'o042700);
`MEM('o004450, 16'o177400);
`MEM('o004452, 16'o110160);
`MEM('o004454, 16'o021660);
`MEM('o004456, 16'o016565);
`MEM('o004460, 16'o177772);
`MEM('o004462, 16'o177770);
`MEM('o004464, 16'o000167);
`MEM('o004466, 16'o000632);
`MEM('o004470, 16'o117500);
`MEM('o004472, 16'o177770);
`MEM('o004474, 16'o120027);
`MEM('o004476, 16'o000042);
`MEM('o004500, 16'o001405);
`MEM('o004502, 16'o117500);
`MEM('o004504, 16'o177770);
`MEM('o004506, 16'o120027);
`MEM('o004510, 16'o000047);
`MEM('o004512, 16'o001155);
`MEM('o004514, 16'o016500);
`MEM('o004516, 16'o177770);
`MEM('o004520, 16'o010001);
`MEM('o004522, 16'o005201);
`MEM('o004524, 16'o010165);
`MEM('o004526, 16'o177770);
`MEM('o004530, 16'o111065);
`MEM('o004532, 16'o177765);
`MEM('o004534, 16'o016565);
`MEM('o004536, 16'o177770);
`MEM('o004540, 16'o177772);
`MEM('o004542, 16'o105065);
`MEM('o004544, 16'o177777);
`MEM('o004546, 16'o000410);
`MEM('o004550, 16'o005265);
`MEM('o004552, 16'o177772);
`MEM('o004554, 16'o116500);
`MEM('o004556, 16'o177777);
`MEM('o004560, 16'o110002);
`MEM('o004562, 16'o105202);
`MEM('o004564, 16'o110265);
`MEM('o004566, 16'o177777);
`MEM('o004570, 16'o117500);
`MEM('o004572, 16'o177772);
`MEM('o004574, 16'o126500);
`MEM('o004576, 16'o177765);
`MEM('o004600, 16'o001411);
`MEM('o004602, 16'o117500);
`MEM('o004604, 16'o177772);
`MEM('o004606, 16'o110046);
`MEM('o004610, 16'o004767);
`MEM('o004612, 16'o174520);
`MEM('o004614, 16'o062706);
`MEM('o004616, 16'o000002);
`MEM('o004620, 16'o105700);
`MEM('o004622, 16'o001352);
`MEM('o004624, 16'o005000);
`MEM('o004626, 16'o156500);
`MEM('o004630, 16'o177776);
`MEM('o004632, 16'o005001);
`MEM('o004634, 16'o156501);
`MEM('o004636, 16'o177777);
`MEM('o004640, 16'o012702);
`MEM('o004642, 16'o000117);
`MEM('o004644, 16'o160102);
`MEM('o004646, 16'o020002);
`MEM('o004650, 16'o002406);
`MEM('o004652, 16'o112767);
`MEM('o004654, 16'o000004);
`MEM('o004656, 16'o013770);
`MEM('o004660, 16'o105000);
`MEM('o004662, 16'o000167);
`MEM('o004664, 16'o000502);
`MEM('o004666, 16'o116500);
`MEM('o004670, 16'o177776);
`MEM('o004672, 16'o110001);
`MEM('o004674, 16'o105201);
`MEM('o004676, 16'o110165);
`MEM('o004700, 16'o177776);
`MEM('o004702, 16'o042700);
`MEM('o004704, 16'o177400);
`MEM('o004706, 16'o112760);
`MEM('o004710, 16'o000044);
`MEM('o004712, 16'o021660);
`MEM('o004714, 16'o116500);
`MEM('o004716, 16'o177776);
`MEM('o004720, 16'o110002);
`MEM('o004722, 16'o105202);
`MEM('o004724, 16'o110265);
`MEM('o004726, 16'o177776);
`MEM('o004730, 16'o042700);
`MEM('o004732, 16'o177400);
`MEM('o004734, 16'o116560);
`MEM('o004736, 16'o177777);
`MEM('o004740, 16'o021660);
`MEM('o004742, 16'o000421);
`MEM('o004744, 16'o016500);
`MEM('o004746, 16'o177770);
`MEM('o004750, 16'o010001);
`MEM('o004752, 16'o005201);
`MEM('o004754, 16'o010165);
`MEM('o004756, 16'o177770);
`MEM('o004760, 16'o111001);
`MEM('o004762, 16'o116500);
`MEM('o004764, 16'o177776);
`MEM('o004766, 16'o110002);
`MEM('o004770, 16'o105202);
`MEM('o004772, 16'o110265);
`MEM('o004774, 16'o177776);
`MEM('o004776, 16'o042700);
`MEM('o005000, 16'o177400);
`MEM('o005002, 16'o110160);
`MEM('o005004, 16'o021660);
`MEM('o005006, 16'o116500);
`MEM('o005010, 16'o177777);
`MEM('o005012, 16'o110001);
`MEM('o005014, 16'o105301);
`MEM('o005016, 16'o110165);
`MEM('o005020, 16'o177777);
`MEM('o005022, 16'o105700);
`MEM('o005024, 16'o001347);
`MEM('o005026, 16'o117500);
`MEM('o005030, 16'o177770);
`MEM('o005032, 16'o126500);
`MEM('o005034, 16'o177765);
`MEM('o005036, 16'o001131);
`MEM('o005040, 16'o005265);
`MEM('o005042, 16'o177770);
`MEM('o005044, 16'o000526);
`MEM('o005046, 16'o117500);
`MEM('o005050, 16'o177772);
`MEM('o005052, 16'o110046);
`MEM('o005054, 16'o004767);
`MEM('o005056, 16'o174424);
`MEM('o005060, 16'o062706);
`MEM('o005062, 16'o000002);
`MEM('o005064, 16'o105700);
`MEM('o005066, 16'o001510);
`MEM('o005070, 16'o126527);
`MEM('o005072, 16'o177776);
`MEM('o005074, 16'o000115);
`MEM('o005076, 16'o101405);
`MEM('o005100, 16'o112767);
`MEM('o005102, 16'o000004);
`MEM('o005104, 16'o013542);
`MEM('o005106, 16'o105000);
`MEM('o005110, 16'o000527);
`MEM('o005112, 16'o126527);
`MEM('o005114, 16'o177776);
`MEM('o005116, 16'o000003);
`MEM('o005120, 16'o101431);
`MEM('o005122, 16'o005000);
`MEM('o005124, 16'o156500);
`MEM('o005126, 16'o177776);
`MEM('o005130, 16'o062700);
`MEM('o005132, 16'o177776);
`MEM('o005134, 16'o116000);
`MEM('o005136, 16'o021660);
`MEM('o005140, 16'o120027);
`MEM('o005142, 16'o000043);
`MEM('o005144, 16'o001017);
`MEM('o005146, 16'o005000);
`MEM('o005150, 16'o156500);
`MEM('o005152, 16'o177776);
`MEM('o005154, 16'o062700);
`MEM('o005156, 16'o177774);
`MEM('o005160, 16'o116000);
`MEM('o005162, 16'o021660);
`MEM('o005164, 16'o120027);
`MEM('o005166, 16'o000043);
`MEM('o005170, 16'o001005);
`MEM('o005172, 16'o112767);
`MEM('o005174, 16'o000024);
`MEM('o005176, 16'o013450);
`MEM('o005200, 16'o105000);
`MEM('o005202, 16'o000472);
`MEM('o005204, 16'o116500);
`MEM('o005206, 16'o177776);
`MEM('o005210, 16'o110002);
`MEM('o005212, 16'o105202);
`MEM('o005214, 16'o110265);
`MEM('o005216, 16'o177776);
`MEM('o005220, 16'o042700);
`MEM('o005222, 16'o177400);
`MEM('o005224, 16'o112760);
`MEM('o005226, 16'o000043);
`MEM('o005230, 16'o021660);
`MEM('o005232, 16'o117500);
`MEM('o005234, 16'o177772);
`MEM('o005236, 16'o110046);
`MEM('o005240, 16'o004767);
`MEM('o005242, 16'o174022);
`MEM('o005244, 16'o062706);
`MEM('o005246, 16'o000002);
`MEM('o005250, 16'o110001);
`MEM('o005252, 16'o116500);
`MEM('o005254, 16'o177776);
`MEM('o005256, 16'o110002);
`MEM('o005260, 16'o105202);
`MEM('o005262, 16'o110265);
`MEM('o005264, 16'o177776);
`MEM('o005266, 16'o042700);
`MEM('o005270, 16'o177400);
`MEM('o005272, 16'o062701);
`MEM('o005274, 16'o177677);
`MEM('o005276, 16'o110160);
`MEM('o005300, 16'o021660);
`MEM('o005302, 16'o005265);
`MEM('o005304, 16'o177770);
`MEM('o005306, 16'o000405);
`MEM('o005310, 16'o112767);
`MEM('o005312, 16'o000024);
`MEM('o005314, 16'o013332);
`MEM('o005316, 16'o105000);
`MEM('o005320, 16'o000423);
`MEM('o005322, 16'o117500);
`MEM('o005324, 16'o177770);
`MEM('o005326, 16'o105700);
`MEM('o005330, 16'o001402);
`MEM('o005332, 16'o000167);
`MEM('o005334, 16'o176020);
`MEM('o005336, 16'o116500);
`MEM('o005340, 16'o177776);
`MEM('o005342, 16'o110001);
`MEM('o005344, 16'o105201);
`MEM('o005346, 16'o110165);
`MEM('o005350, 16'o177776);
`MEM('o005352, 16'o042700);
`MEM('o005354, 16'o177400);
`MEM('o005356, 16'o112760);
`MEM('o005360, 16'o000045);
`MEM('o005362, 16'o021660);
`MEM('o005364, 16'o116500);
`MEM('o005366, 16'o177776);
`MEM('o005370, 16'o010506);
`MEM('o005372, 16'o012605);
`MEM('o005374, 16'o012602);
`MEM('o005376, 16'o000207);
`MEM('o005400, 16'o010546);
`MEM('o005402, 16'o010605);
`MEM('o005404, 16'o062706);
`MEM('o005406, 16'o177776);
`MEM('o005410, 16'o012765);
`MEM('o005412, 16'o022164);
`MEM('o005414, 16'o177776);
`MEM('o005416, 16'o000406);
`MEM('o005420, 16'o117500);
`MEM('o005422, 16'o177776);
`MEM('o005424, 16'o042700);
`MEM('o005426, 16'o177400);
`MEM('o005430, 16'o060065);
`MEM('o005432, 16'o177776);
`MEM('o005434, 16'o117500);
`MEM('o005436, 16'o177776);
`MEM('o005440, 16'o105700);
`MEM('o005442, 16'o001366);
`MEM('o005444, 16'o012700);
`MEM('o005446, 16'o024164);
`MEM('o005450, 16'o166500);
`MEM('o005452, 16'o177776);
`MEM('o005454, 16'o005300);
`MEM('o005456, 16'o010506);
`MEM('o005460, 16'o012605);
`MEM('o005462, 16'o000207);
`MEM('o005464, 16'o010546);
`MEM('o005466, 16'o010605);
`MEM('o005470, 16'o117500);
`MEM('o005472, 16'o000004);
`MEM('o005474, 16'o105700);
`MEM('o005476, 16'o001003);
`MEM('o005500, 16'o012700);
`MEM('o005502, 16'o077777);
`MEM('o005504, 16'o000420);
`MEM('o005506, 16'o016500);
`MEM('o005510, 16'o000004);
`MEM('o005512, 16'o005200);
`MEM('o005514, 16'o111000);
`MEM('o005516, 16'o005001);
`MEM('o005520, 16'o150001);
`MEM('o005522, 16'o016500);
`MEM('o005524, 16'o000004);
`MEM('o005526, 16'o062700);
`MEM('o005530, 16'o000002);
`MEM('o005532, 16'o111000);
`MEM('o005534, 16'o042700);
`MEM('o005536, 16'o177400);
`MEM('o005540, 16'o072027);
`MEM('o005542, 16'o000010);
`MEM('o005544, 16'o050100);
`MEM('o005546, 16'o012605);
`MEM('o005550, 16'o000207);
`MEM('o005552, 16'o010546);
`MEM('o005554, 16'o010605);
`MEM('o005556, 16'o062706);
`MEM('o005560, 16'o177776);
`MEM('o005562, 16'o012765);
`MEM('o005564, 16'o022164);
`MEM('o005566, 16'o177776);
`MEM('o005570, 16'o000417);
`MEM('o005572, 16'o016546);
`MEM('o005574, 16'o177776);
`MEM('o005576, 16'o004767);
`MEM('o005600, 16'o177662);
`MEM('o005602, 16'o062706);
`MEM('o005604, 16'o000002);
`MEM('o005606, 16'o026500);
`MEM('o005610, 16'o000004);
`MEM('o005612, 16'o003413);
`MEM('o005614, 16'o117500);
`MEM('o005616, 16'o177776);
`MEM('o005620, 16'o042700);
`MEM('o005622, 16'o177400);
`MEM('o005624, 16'o060065);
`MEM('o005626, 16'o177776);
`MEM('o005630, 16'o117500);
`MEM('o005632, 16'o177776);
`MEM('o005634, 16'o105700);
`MEM('o005636, 16'o001355);
`MEM('o005640, 16'o000401);
`MEM('o005642, 16'o000240);
`MEM('o005644, 16'o016500);
`MEM('o005646, 16'o177776);
`MEM('o005650, 16'o010506);
`MEM('o005652, 16'o012605);
`MEM('o005654, 16'o000207);
`MEM('o005656, 16'o010246);
`MEM('o005660, 16'o010546);
`MEM('o005662, 16'o010605);
`MEM('o005664, 16'o062706);
`MEM('o005666, 16'o177770);
`MEM('o005670, 16'o004767);
`MEM('o005672, 16'o177504);
`MEM('o005674, 16'o116701);
`MEM('o005676, 16'o013760);
`MEM('o005700, 16'o042701);
`MEM('o005702, 16'o177400);
`MEM('o005704, 16'o020001);
`MEM('o005706, 16'o002005);
`MEM('o005710, 16'o112767);
`MEM('o005712, 16'o000005);
`MEM('o005714, 16'o012732);
`MEM('o005716, 16'o000167);
`MEM('o005720, 16'o000524);
`MEM('o005722, 16'o012746);
`MEM('o005724, 16'o021660);
`MEM('o005726, 16'o004767);
`MEM('o005730, 16'o177532);
`MEM('o005732, 16'o062706);
`MEM('o005734, 16'o000002);
`MEM('o005736, 16'o010046);
`MEM('o005740, 16'o004767);
`MEM('o005742, 16'o177606);
`MEM('o005744, 16'o062706);
`MEM('o005746, 16'o000002);
`MEM('o005750, 16'o010065);
`MEM('o005752, 16'o177770);
`MEM('o005754, 16'o016546);
`MEM('o005756, 16'o177770);
`MEM('o005760, 16'o004767);
`MEM('o005762, 16'o177500);
`MEM('o005764, 16'o062706);
`MEM('o005766, 16'o000002);
`MEM('o005770, 16'o010002);
`MEM('o005772, 16'o012746);
`MEM('o005774, 16'o021660);
`MEM('o005776, 16'o004767);
`MEM('o006000, 16'o177462);
`MEM('o006002, 16'o062706);
`MEM('o006004, 16'o000002);
`MEM('o006006, 16'o020200);
`MEM('o006010, 16'o001056);
`MEM('o006012, 16'o016565);
`MEM('o006014, 16'o177770);
`MEM('o006016, 16'o177776);
`MEM('o006020, 16'o117500);
`MEM('o006022, 16'o177776);
`MEM('o006024, 16'o042700);
`MEM('o006026, 16'o177400);
`MEM('o006030, 16'o016501);
`MEM('o006032, 16'o177776);
`MEM('o006034, 16'o060001);
`MEM('o006036, 16'o010165);
`MEM('o006040, 16'o177774);
`MEM('o006042, 16'o000426);
`MEM('o006044, 16'o016501);
`MEM('o006046, 16'o177774);
`MEM('o006050, 16'o010102);
`MEM('o006052, 16'o005202);
`MEM('o006054, 16'o010265);
`MEM('o006056, 16'o177774);
`MEM('o006060, 16'o016500);
`MEM('o006062, 16'o177776);
`MEM('o006064, 16'o010002);
`MEM('o006066, 16'o005202);
`MEM('o006070, 16'o010265);
`MEM('o006072, 16'o177776);
`MEM('o006074, 16'o111101);
`MEM('o006076, 16'o110110);
`MEM('o006100, 16'o016500);
`MEM('o006102, 16'o177772);
`MEM('o006104, 16'o010001);
`MEM('o006106, 16'o005301);
`MEM('o006110, 16'o010165);
`MEM('o006112, 16'o177772);
`MEM('o006114, 16'o005700);
`MEM('o006116, 16'o001352);
`MEM('o006120, 16'o117500);
`MEM('o006122, 16'o177774);
`MEM('o006124, 16'o005001);
`MEM('o006126, 16'o150001);
`MEM('o006130, 16'o010165);
`MEM('o006132, 16'o177772);
`MEM('o006134, 16'o005765);
`MEM('o006136, 16'o177772);
`MEM('o006140, 16'o001357);
`MEM('o006142, 16'o105075);
`MEM('o006144, 16'o177776);
`MEM('o006146, 16'o116700);
`MEM('o006150, 16'o013506);
`MEM('o006152, 16'o120027);
`MEM('o006154, 16'o000004);
`MEM('o006156, 16'o001532);
`MEM('o006160, 16'o016565);
`MEM('o006162, 16'o177770);
`MEM('o006164, 16'o177776);
`MEM('o006166, 16'o000406);
`MEM('o006170, 16'o117500);
`MEM('o006172, 16'o177776);
`MEM('o006174, 16'o042700);
`MEM('o006176, 16'o177400);
`MEM('o006200, 16'o060065);
`MEM('o006202, 16'o177776);
`MEM('o006204, 16'o117500);
`MEM('o006206, 16'o177776);
`MEM('o006210, 16'o105700);
`MEM('o006212, 16'o001366);
`MEM('o006214, 16'o016500);
`MEM('o006216, 16'o177776);
`MEM('o006220, 16'o166500);
`MEM('o006222, 16'o177770);
`MEM('o006224, 16'o010002);
`MEM('o006226, 16'o005202);
`MEM('o006230, 16'o010265);
`MEM('o006232, 16'o177772);
`MEM('o006234, 16'o116700);
`MEM('o006236, 16'o013420);
`MEM('o006240, 16'o042700);
`MEM('o006242, 16'o177400);
`MEM('o006244, 16'o016501);
`MEM('o006246, 16'o177776);
`MEM('o006250, 16'o060001);
`MEM('o006252, 16'o010165);
`MEM('o006254, 16'o177774);
`MEM('o006256, 16'o000416);
`MEM('o006260, 16'o016501);
`MEM('o006262, 16'o177776);
`MEM('o006264, 16'o010102);
`MEM('o006266, 16'o005302);
`MEM('o006270, 16'o010265);
`MEM('o006272, 16'o177776);
`MEM('o006274, 16'o016500);
`MEM('o006276, 16'o177774);
`MEM('o006300, 16'o010002);
`MEM('o006302, 16'o005302);
`MEM('o006304, 16'o010265);
`MEM('o006306, 16'o177774);
`MEM('o006310, 16'o111101);
`MEM('o006312, 16'o110110);
`MEM('o006314, 16'o016500);
`MEM('o006316, 16'o177772);
`MEM('o006320, 16'o010001);
`MEM('o006322, 16'o005301);
`MEM('o006324, 16'o010165);
`MEM('o006326, 16'o177772);
`MEM('o006330, 16'o005700);
`MEM('o006332, 16'o001352);
`MEM('o006334, 16'o116700);
`MEM('o006336, 16'o013320);
`MEM('o006340, 16'o005001);
`MEM('o006342, 16'o150001);
`MEM('o006344, 16'o010165);
`MEM('o006346, 16'o177772);
`MEM('o006350, 16'o016565);
`MEM('o006352, 16'o177770);
`MEM('o006354, 16'o177776);
`MEM('o006356, 16'o012765);
`MEM('o006360, 16'o021660);
`MEM('o006362, 16'o177774);
`MEM('o006364, 16'o000416);
`MEM('o006366, 16'o016501);
`MEM('o006370, 16'o177774);
`MEM('o006372, 16'o010102);
`MEM('o006374, 16'o005202);
`MEM('o006376, 16'o010265);
`MEM('o006400, 16'o177774);
`MEM('o006402, 16'o016500);
`MEM('o006404, 16'o177776);
`MEM('o006406, 16'o010002);
`MEM('o006410, 16'o005202);
`MEM('o006412, 16'o010265);
`MEM('o006414, 16'o177776);
`MEM('o006416, 16'o111101);
`MEM('o006420, 16'o110110);
`MEM('o006422, 16'o016500);
`MEM('o006424, 16'o177772);
`MEM('o006426, 16'o010001);
`MEM('o006430, 16'o005301);
`MEM('o006432, 16'o010165);
`MEM('o006434, 16'o177772);
`MEM('o006436, 16'o005700);
`MEM('o006440, 16'o001352);
`MEM('o006442, 16'o000401);
`MEM('o006444, 16'o000240);
`MEM('o006446, 16'o010506);
`MEM('o006450, 16'o012605);
`MEM('o006452, 16'o012602);
`MEM('o006454, 16'o000207);
`MEM('o006456, 16'o010546);
`MEM('o006460, 16'o010605);
`MEM('o006462, 16'o062706);
`MEM('o006464, 16'o177776);
`MEM('o006466, 16'o000167);
`MEM('o006470, 16'o001042);
`MEM('o006472, 16'o117500);
`MEM('o006474, 16'o000004);
`MEM('o006476, 16'o120027);
`MEM('o006500, 16'o000041);
`MEM('o006502, 16'o101114);
`MEM('o006504, 16'o117500);
`MEM('o006506, 16'o000004);
`MEM('o006510, 16'o042700);
`MEM('o006512, 16'o177400);
`MEM('o006514, 16'o006300);
`MEM('o006516, 16'o062700);
`MEM('o006520, 16'o020502);
`MEM('o006522, 16'o011000);
`MEM('o006524, 16'o010046);
`MEM('o006526, 16'o004767);
`MEM('o006530, 16'o173032);
`MEM('o006532, 16'o062706);
`MEM('o006534, 16'o000002);
`MEM('o006536, 16'o117500);
`MEM('o006540, 16'o000004);
`MEM('o006542, 16'o112746);
`MEM('o006544, 16'o000023);
`MEM('o006546, 16'o012746);
`MEM('o006550, 16'o020606);
`MEM('o006552, 16'o110046);
`MEM('o006554, 16'o004767);
`MEM('o006556, 16'o172422);
`MEM('o006560, 16'o062706);
`MEM('o006562, 16'o000006);
`MEM('o006564, 16'o105700);
`MEM('o006566, 16'o001006);
`MEM('o006570, 16'o012746);
`MEM('o006572, 16'o000040);
`MEM('o006574, 16'o004767);
`MEM('o006576, 16'o172210);
`MEM('o006600, 16'o062706);
`MEM('o006602, 16'o000002);
`MEM('o006604, 16'o117500);
`MEM('o006606, 16'o000004);
`MEM('o006610, 16'o120027);
`MEM('o006612, 16'o000010);
`MEM('o006614, 16'o001043);
`MEM('o006616, 16'o005265);
`MEM('o006620, 16'o000004);
`MEM('o006622, 16'o016500);
`MEM('o006624, 16'o000004);
`MEM('o006626, 16'o010001);
`MEM('o006630, 16'o005201);
`MEM('o006632, 16'o010165);
`MEM('o006634, 16'o000004);
`MEM('o006636, 16'o111065);
`MEM('o006640, 16'o177777);
`MEM('o006642, 16'o000416);
`MEM('o006644, 16'o016500);
`MEM('o006646, 16'o000004);
`MEM('o006650, 16'o010001);
`MEM('o006652, 16'o005201);
`MEM('o006654, 16'o010165);
`MEM('o006656, 16'o000004);
`MEM('o006660, 16'o111000);
`MEM('o006662, 16'o042700);
`MEM('o006664, 16'o177400);
`MEM('o006666, 16'o010046);
`MEM('o006670, 16'o004767);
`MEM('o006672, 16'o172114);
`MEM('o006674, 16'o062706);
`MEM('o006676, 16'o000002);
`MEM('o006700, 16'o116500);
`MEM('o006702, 16'o177777);
`MEM('o006704, 16'o110001);
`MEM('o006706, 16'o105301);
`MEM('o006710, 16'o110165);
`MEM('o006712, 16'o177777);
`MEM('o006714, 16'o105700);
`MEM('o006716, 16'o001352);
`MEM('o006720, 16'o000167);
`MEM('o006722, 16'o000626);
`MEM('o006724, 16'o005265);
`MEM('o006726, 16'o000004);
`MEM('o006730, 16'o000167);
`MEM('o006732, 16'o000600);
`MEM('o006734, 16'o117500);
`MEM('o006736, 16'o000004);
`MEM('o006740, 16'o120027);
`MEM('o006742, 16'o000042);
`MEM('o006744, 16'o001057);
`MEM('o006746, 16'o005265);
`MEM('o006750, 16'o000004);
`MEM('o006752, 16'o117500);
`MEM('o006754, 16'o000004);
`MEM('o006756, 16'o005001);
`MEM('o006760, 16'o150001);
`MEM('o006762, 16'o016500);
`MEM('o006764, 16'o000004);
`MEM('o006766, 16'o005200);
`MEM('o006770, 16'o111000);
`MEM('o006772, 16'o042700);
`MEM('o006774, 16'o177400);
`MEM('o006776, 16'o072027);
`MEM('o007000, 16'o000010);
`MEM('o007002, 16'o050100);
`MEM('o007004, 16'o005046);
`MEM('o007006, 16'o010046);
`MEM('o007010, 16'o004767);
`MEM('o007012, 16'o173220);
`MEM('o007014, 16'o062706);
`MEM('o007016, 16'o000004);
`MEM('o007020, 16'o062765);
`MEM('o007022, 16'o000002);
`MEM('o007024, 16'o000004);
`MEM('o007026, 16'o117500);
`MEM('o007030, 16'o000004);
`MEM('o007032, 16'o112746);
`MEM('o007034, 16'o000017);
`MEM('o007036, 16'o012746);
`MEM('o007040, 16'o020631);
`MEM('o007042, 16'o110046);
`MEM('o007044, 16'o004767);
`MEM('o007046, 16'o172132);
`MEM('o007050, 16'o062706);
`MEM('o007052, 16'o000006);
`MEM('o007054, 16'o105700);
`MEM('o007056, 16'o001402);
`MEM('o007060, 16'o000167);
`MEM('o007062, 16'o000450);
`MEM('o007064, 16'o012746);
`MEM('o007066, 16'o000040);
`MEM('o007070, 16'o004767);
`MEM('o007072, 16'o171714);
`MEM('o007074, 16'o062706);
`MEM('o007076, 16'o000002);
`MEM('o007100, 16'o000167);
`MEM('o007102, 16'o000430);
`MEM('o007104, 16'o117500);
`MEM('o007106, 16'o000004);
`MEM('o007110, 16'o120027);
`MEM('o007112, 16'o000043);
`MEM('o007114, 16'o001046);
`MEM('o007116, 16'o005265);
`MEM('o007120, 16'o000004);
`MEM('o007122, 16'o016500);
`MEM('o007124, 16'o000004);
`MEM('o007126, 16'o010001);
`MEM('o007130, 16'o005201);
`MEM('o007132, 16'o010165);
`MEM('o007134, 16'o000004);
`MEM('o007136, 16'o111000);
`MEM('o007140, 16'o042700);
`MEM('o007142, 16'o177400);
`MEM('o007144, 16'o062700);
`MEM('o007146, 16'o000101);
`MEM('o007150, 16'o010046);
`MEM('o007152, 16'o004767);
`MEM('o007154, 16'o171632);
`MEM('o007156, 16'o062706);
`MEM('o007160, 16'o000002);
`MEM('o007162, 16'o117500);
`MEM('o007164, 16'o000004);
`MEM('o007166, 16'o112746);
`MEM('o007170, 16'o000017);
`MEM('o007172, 16'o012746);
`MEM('o007174, 16'o020631);
`MEM('o007176, 16'o110046);
`MEM('o007200, 16'o004767);
`MEM('o007202, 16'o171776);
`MEM('o007204, 16'o062706);
`MEM('o007206, 16'o000006);
`MEM('o007210, 16'o105700);
`MEM('o007212, 16'o001150);
`MEM('o007214, 16'o012746);
`MEM('o007216, 16'o000040);
`MEM('o007220, 16'o004767);
`MEM('o007222, 16'o171564);
`MEM('o007224, 16'o062706);
`MEM('o007226, 16'o000002);
`MEM('o007230, 16'o000541);
`MEM('o007232, 16'o117500);
`MEM('o007234, 16'o000004);
`MEM('o007236, 16'o120027);
`MEM('o007240, 16'o000044);
`MEM('o007242, 16'o001130);
`MEM('o007244, 16'o112765);
`MEM('o007246, 16'o000042);
`MEM('o007250, 16'o177776);
`MEM('o007252, 16'o005265);
`MEM('o007254, 16'o000004);
`MEM('o007256, 16'o117565);
`MEM('o007260, 16'o000004);
`MEM('o007262, 16'o177777);
`MEM('o007264, 16'o000423);
`MEM('o007266, 16'o005000);
`MEM('o007270, 16'o156500);
`MEM('o007272, 16'o177777);
`MEM('o007274, 16'o066500);
`MEM('o007276, 16'o000004);
`MEM('o007300, 16'o111000);
`MEM('o007302, 16'o120027);
`MEM('o007304, 16'o000042);
`MEM('o007306, 16'o001004);
`MEM('o007310, 16'o112765);
`MEM('o007312, 16'o000047);
`MEM('o007314, 16'o177776);
`MEM('o007316, 16'o000411);
`MEM('o007320, 16'o116500);
`MEM('o007322, 16'o177777);
`MEM('o007324, 16'o110001);
`MEM('o007326, 16'o105301);
`MEM('o007330, 16'o110165);
`MEM('o007332, 16'o177777);
`MEM('o007334, 16'o105765);
`MEM('o007336, 16'o177777);
`MEM('o007340, 16'o001352);
`MEM('o007342, 16'o116500);
`MEM('o007344, 16'o177776);
`MEM('o007346, 16'o010046);
`MEM('o007350, 16'o004767);
`MEM('o007352, 16'o171434);
`MEM('o007354, 16'o062706);
`MEM('o007356, 16'o000002);
`MEM('o007360, 16'o016500);
`MEM('o007362, 16'o000004);
`MEM('o007364, 16'o010001);
`MEM('o007366, 16'o005201);
`MEM('o007370, 16'o010165);
`MEM('o007372, 16'o000004);
`MEM('o007374, 16'o111065);
`MEM('o007376, 16'o177777);
`MEM('o007400, 16'o000416);
`MEM('o007402, 16'o016500);
`MEM('o007404, 16'o000004);
`MEM('o007406, 16'o010001);
`MEM('o007410, 16'o005201);
`MEM('o007412, 16'o010165);
`MEM('o007414, 16'o000004);
`MEM('o007416, 16'o111000);
`MEM('o007420, 16'o042700);
`MEM('o007422, 16'o177400);
`MEM('o007424, 16'o010046);
`MEM('o007426, 16'o004767);
`MEM('o007430, 16'o171356);
`MEM('o007432, 16'o062706);
`MEM('o007434, 16'o000002);
`MEM('o007436, 16'o116500);
`MEM('o007440, 16'o177777);
`MEM('o007442, 16'o110001);
`MEM('o007444, 16'o105301);
`MEM('o007446, 16'o110165);
`MEM('o007450, 16'o177777);
`MEM('o007452, 16'o105700);
`MEM('o007454, 16'o001352);
`MEM('o007456, 16'o116500);
`MEM('o007460, 16'o177776);
`MEM('o007462, 16'o010046);
`MEM('o007464, 16'o004767);
`MEM('o007466, 16'o171320);
`MEM('o007470, 16'o062706);
`MEM('o007472, 16'o000002);
`MEM('o007474, 16'o117500);
`MEM('o007476, 16'o000004);
`MEM('o007500, 16'o120027);
`MEM('o007502, 16'o000043);
`MEM('o007504, 16'o001013);
`MEM('o007506, 16'o012746);
`MEM('o007510, 16'o000040);
`MEM('o007512, 16'o004767);
`MEM('o007514, 16'o171272);
`MEM('o007516, 16'o062706);
`MEM('o007520, 16'o000002);
`MEM('o007522, 16'o000404);
`MEM('o007524, 16'o112767);
`MEM('o007526, 16'o000025);
`MEM('o007530, 16'o011116);
`MEM('o007532, 16'o000407);
`MEM('o007534, 16'o117500);
`MEM('o007536, 16'o000004);
`MEM('o007540, 16'o120027);
`MEM('o007542, 16'o000045);
`MEM('o007544, 16'o001402);
`MEM('o007546, 16'o000167);
`MEM('o007550, 16'o176720);
`MEM('o007552, 16'o010506);
`MEM('o007554, 16'o012605);
`MEM('o007556, 16'o000207);
`MEM('o007560, 16'o010546);
`MEM('o007562, 16'o010605);
`MEM('o007564, 16'o062706);
`MEM('o007566, 16'o177776);
`MEM('o007570, 16'o016700);
`MEM('o007572, 16'o014372);
`MEM('o007574, 16'o111000);
`MEM('o007576, 16'o120027);
`MEM('o007600, 16'o000023);
`MEM('o007602, 16'o001405);
`MEM('o007604, 16'o112767);
`MEM('o007606, 16'o000021);
`MEM('o007610, 16'o011036);
`MEM('o007612, 16'o005000);
`MEM('o007614, 16'o000441);
`MEM('o007616, 16'o016700);
`MEM('o007620, 16'o014344);
`MEM('o007622, 16'o005200);
`MEM('o007624, 16'o010067);
`MEM('o007626, 16'o014336);
`MEM('o007630, 16'o004767);
`MEM('o007632, 16'o001326);
`MEM('o007634, 16'o010065);
`MEM('o007636, 16'o177776);
`MEM('o007640, 16'o116700);
`MEM('o007642, 16'o011004);
`MEM('o007644, 16'o105700);
`MEM('o007646, 16'o001402);
`MEM('o007650, 16'o005000);
`MEM('o007652, 16'o000422);
`MEM('o007654, 16'o016700);
`MEM('o007656, 16'o014306);
`MEM('o007660, 16'o111000);
`MEM('o007662, 16'o120027);
`MEM('o007664, 16'o000024);
`MEM('o007666, 16'o001405);
`MEM('o007670, 16'o112767);
`MEM('o007672, 16'o000021);
`MEM('o007674, 16'o010752);
`MEM('o007676, 16'o005000);
`MEM('o007700, 16'o000407);
`MEM('o007702, 16'o016700);
`MEM('o007704, 16'o014260);
`MEM('o007706, 16'o005200);
`MEM('o007710, 16'o010067);
`MEM('o007712, 16'o014252);
`MEM('o007714, 16'o016500);
`MEM('o007716, 16'o177776);
`MEM('o007720, 16'o010506);
`MEM('o007722, 16'o012605);
`MEM('o007724, 16'o000207);
`MEM('o007726, 16'o010246);
`MEM('o007730, 16'o010546);
`MEM('o007732, 16'o010605);
`MEM('o007734, 16'o062706);
`MEM('o007736, 16'o177776);
`MEM('o007740, 16'o016700);
`MEM('o007742, 16'o014222);
`MEM('o007744, 16'o111000);
`MEM('o007746, 16'o042700);
`MEM('o007750, 16'o177400);
`MEM('o007752, 16'o062700);
`MEM('o007754, 16'o177761);
`MEM('o007756, 16'o020027);
`MEM('o007760, 16'o000024);
`MEM('o007762, 16'o101402);
`MEM('o007764, 16'o000167);
`MEM('o007766, 16'o000512);
`MEM('o007770, 16'o006300);
`MEM('o007772, 16'o062700);
`MEM('o007774, 16'o024246);
`MEM('o007776, 16'o011000);
`MEM('o010000, 16'o000110);
`MEM('o010002, 16'o016700);
`MEM('o010004, 16'o014160);
`MEM('o010006, 16'o005200);
`MEM('o010010, 16'o010067);
`MEM('o010012, 16'o014152);
`MEM('o010014, 16'o016700);
`MEM('o010016, 16'o014146);
`MEM('o010020, 16'o111000);
`MEM('o010022, 16'o005001);
`MEM('o010024, 16'o150001);
`MEM('o010026, 16'o016700);
`MEM('o010030, 16'o014134);
`MEM('o010032, 16'o005200);
`MEM('o010034, 16'o111000);
`MEM('o010036, 16'o042700);
`MEM('o010040, 16'o177400);
`MEM('o010042, 16'o072027);
`MEM('o010044, 16'o000010);
`MEM('o010046, 16'o010102);
`MEM('o010050, 16'o050002);
`MEM('o010052, 16'o010265);
`MEM('o010054, 16'o177776);
`MEM('o010056, 16'o016700);
`MEM('o010060, 16'o014104);
`MEM('o010062, 16'o062700);
`MEM('o010064, 16'o000002);
`MEM('o010066, 16'o010067);
`MEM('o010070, 16'o014074);
`MEM('o010072, 16'o000167);
`MEM('o010074, 16'o000426);
`MEM('o010076, 16'o016700);
`MEM('o010100, 16'o014064);
`MEM('o010102, 16'o005200);
`MEM('o010104, 16'o010067);
`MEM('o010106, 16'o014056);
`MEM('o010110, 16'o004767);
`MEM('o010112, 16'o177612);
`MEM('o010114, 16'o010065);
`MEM('o010116, 16'o177776);
`MEM('o010120, 16'o000167);
`MEM('o010122, 16'o000400);
`MEM('o010124, 16'o016700);
`MEM('o010126, 16'o014036);
`MEM('o010130, 16'o005200);
`MEM('o010132, 16'o010067);
`MEM('o010134, 16'o014030);
`MEM('o010136, 16'o004767);
`MEM('o010140, 16'o177564);
`MEM('o010142, 16'o010001);
`MEM('o010144, 16'o005401);
`MEM('o010146, 16'o010165);
`MEM('o010150, 16'o177776);
`MEM('o010152, 16'o000167);
`MEM('o010154, 16'o000346);
`MEM('o010156, 16'o016700);
`MEM('o010160, 16'o014004);
`MEM('o010162, 16'o005200);
`MEM('o010164, 16'o010067);
`MEM('o010166, 16'o013776);
`MEM('o010170, 16'o016700);
`MEM('o010172, 16'o013772);
`MEM('o010174, 16'o010001);
`MEM('o010176, 16'o005201);
`MEM('o010200, 16'o010167);
`MEM('o010202, 16'o013762);
`MEM('o010204, 16'o111000);
`MEM('o010206, 16'o042700);
`MEM('o010210, 16'o177400);
`MEM('o010212, 16'o006300);
`MEM('o010214, 16'o062700);
`MEM('o010216, 16'o022000);
`MEM('o010220, 16'o011065);
`MEM('o010222, 16'o177776);
`MEM('o010224, 16'o000537);
`MEM('o010226, 16'o004767);
`MEM('o010230, 16'o177326);
`MEM('o010232, 16'o010065);
`MEM('o010234, 16'o177776);
`MEM('o010236, 16'o000532);
`MEM('o010240, 16'o016700);
`MEM('o010242, 16'o013722);
`MEM('o010244, 16'o005200);
`MEM('o010246, 16'o010067);
`MEM('o010250, 16'o013714);
`MEM('o010252, 16'o004767);
`MEM('o010254, 16'o177302);
`MEM('o010256, 16'o010065);
`MEM('o010260, 16'o177776);
`MEM('o010262, 16'o116700);
`MEM('o010264, 16'o010362);
`MEM('o010266, 16'o105700);
`MEM('o010270, 16'o001110);
`MEM('o010272, 16'o026527);
`MEM('o010274, 16'o177776);
`MEM('o010276, 16'o000037);
`MEM('o010300, 16'o003404);
`MEM('o010302, 16'o112767);
`MEM('o010304, 16'o000003);
`MEM('o010306, 16'o010340);
`MEM('o010310, 16'o000505);
`MEM('o010312, 16'o016500);
`MEM('o010314, 16'o177776);
`MEM('o010316, 16'o006300);
`MEM('o010320, 16'o062700);
`MEM('o010322, 16'o022064);
`MEM('o010324, 16'o011065);
`MEM('o010326, 16'o177776);
`MEM('o010330, 16'o000475);
`MEM('o010332, 16'o016700);
`MEM('o010334, 16'o013630);
`MEM('o010336, 16'o005200);
`MEM('o010340, 16'o010067);
`MEM('o010342, 16'o013622);
`MEM('o010344, 16'o004767);
`MEM('o010346, 16'o177210);
`MEM('o010350, 16'o010065);
`MEM('o010352, 16'o177776);
`MEM('o010354, 16'o116700);
`MEM('o010356, 16'o010270);
`MEM('o010360, 16'o105700);
`MEM('o010362, 16'o001055);
`MEM('o010364, 16'o005765);
`MEM('o010366, 16'o177776);
`MEM('o010370, 16'o002054);
`MEM('o010372, 16'o005465);
`MEM('o010374, 16'o177776);
`MEM('o010376, 16'o000451);
`MEM('o010400, 16'o016700);
`MEM('o010402, 16'o013562);
`MEM('o010404, 16'o005200);
`MEM('o010406, 16'o010067);
`MEM('o010410, 16'o013554);
`MEM('o010412, 16'o016700);
`MEM('o010414, 16'o013550);
`MEM('o010416, 16'o111000);
`MEM('o010420, 16'o120027);
`MEM('o010422, 16'o000023);
`MEM('o010424, 16'o001007);
`MEM('o010426, 16'o016700);
`MEM('o010430, 16'o013534);
`MEM('o010432, 16'o005200);
`MEM('o010434, 16'o111000);
`MEM('o010436, 16'o120027);
`MEM('o010440, 16'o000024);
`MEM('o010442, 16'o001404);
`MEM('o010444, 16'o112767);
`MEM('o010446, 16'o000021);
`MEM('o010450, 16'o010176);
`MEM('o010452, 16'o000424);
`MEM('o010454, 16'o016700);
`MEM('o010456, 16'o013506);
`MEM('o010460, 16'o062700);
`MEM('o010462, 16'o000002);
`MEM('o010464, 16'o010067);
`MEM('o010466, 16'o013476);
`MEM('o010470, 16'o004767);
`MEM('o010472, 16'o174704);
`MEM('o010474, 16'o010065);
`MEM('o010476, 16'o177776);
`MEM('o010500, 16'o000411);
`MEM('o010502, 16'o112767);
`MEM('o010504, 16'o000024);
`MEM('o010506, 16'o010140);
`MEM('o010510, 16'o000405);
`MEM('o010512, 16'o000240);
`MEM('o010514, 16'o000403);
`MEM('o010516, 16'o000240);
`MEM('o010520, 16'o000401);
`MEM('o010522, 16'o000240);
`MEM('o010524, 16'o016500);
`MEM('o010526, 16'o177776);
`MEM('o010530, 16'o010506);
`MEM('o010532, 16'o012605);
`MEM('o010534, 16'o012602);
`MEM('o010536, 16'o000207);
`MEM('o010540, 16'o010546);
`MEM('o010542, 16'o010605);
`MEM('o010544, 16'o062706);
`MEM('o010546, 16'o177774);
`MEM('o010550, 16'o004767);
`MEM('o010552, 16'o177152);
`MEM('o010554, 16'o010065);
`MEM('o010556, 16'o177776);
`MEM('o010560, 16'o116700);
`MEM('o010562, 16'o010064);
`MEM('o010564, 16'o105700);
`MEM('o010566, 16'o001403);
`MEM('o010570, 16'o012700);
`MEM('o010572, 16'o177777);
`MEM('o010574, 16'o000474);
`MEM('o010576, 16'o016700);
`MEM('o010600, 16'o013364);
`MEM('o010602, 16'o111000);
`MEM('o010604, 16'o042700);
`MEM('o010606, 16'o177400);
`MEM('o010610, 16'o020027);
`MEM('o010612, 16'o000021);
`MEM('o010614, 16'o001404);
`MEM('o010616, 16'o020027);
`MEM('o010620, 16'o000022);
`MEM('o010622, 16'o001423);
`MEM('o010624, 16'o000454);
`MEM('o010626, 16'o016700);
`MEM('o010630, 16'o013334);
`MEM('o010632, 16'o005200);
`MEM('o010634, 16'o010067);
`MEM('o010636, 16'o013326);
`MEM('o010640, 16'o004767);
`MEM('o010642, 16'o177062);
`MEM('o010644, 16'o010065);
`MEM('o010646, 16'o177774);
`MEM('o010650, 16'o016500);
`MEM('o010652, 16'o177776);
`MEM('o010654, 16'o016501);
`MEM('o010656, 16'o177774);
`MEM('o010660, 16'o070100);
`MEM('o010662, 16'o010100);
`MEM('o010664, 16'o010065);
`MEM('o010666, 16'o177776);
`MEM('o010670, 16'o000435);
`MEM('o010672, 16'o016700);
`MEM('o010674, 16'o013270);
`MEM('o010676, 16'o005200);
`MEM('o010700, 16'o010067);
`MEM('o010702, 16'o013262);
`MEM('o010704, 16'o004767);
`MEM('o010706, 16'o177016);
`MEM('o010710, 16'o010065);
`MEM('o010712, 16'o177774);
`MEM('o010714, 16'o005765);
`MEM('o010716, 16'o177774);
`MEM('o010720, 16'o001006);
`MEM('o010722, 16'o112767);
`MEM('o010724, 16'o000001);
`MEM('o010726, 16'o007720);
`MEM('o010730, 16'o012700);
`MEM('o010732, 16'o177777);
`MEM('o010734, 16'o000414);
`MEM('o010736, 16'o016501);
`MEM('o010740, 16'o177776);
`MEM('o010742, 16'o006700);
`MEM('o010744, 16'o071065);
`MEM('o010746, 16'o177774);
`MEM('o010750, 16'o010065);
`MEM('o010752, 16'o177776);
`MEM('o010754, 16'o000403);
`MEM('o010756, 16'o016500);
`MEM('o010760, 16'o177776);
`MEM('o010762, 16'o000401);
`MEM('o010764, 16'o000704);
`MEM('o010766, 16'o010506);
`MEM('o010770, 16'o012605);
`MEM('o010772, 16'o000207);
`MEM('o010774, 16'o010546);
`MEM('o010776, 16'o010605);
`MEM('o011000, 16'o062706);
`MEM('o011002, 16'o177774);
`MEM('o011004, 16'o004767);
`MEM('o011006, 16'o177530);
`MEM('o011010, 16'o010065);
`MEM('o011012, 16'o177776);
`MEM('o011014, 16'o116700);
`MEM('o011016, 16'o007630);
`MEM('o011020, 16'o105700);
`MEM('o011022, 16'o001403);
`MEM('o011024, 16'o012700);
`MEM('o011026, 16'o177777);
`MEM('o011030, 16'o000451);
`MEM('o011032, 16'o016700);
`MEM('o011034, 16'o013130);
`MEM('o011036, 16'o111000);
`MEM('o011040, 16'o042700);
`MEM('o011042, 16'o177400);
`MEM('o011044, 16'o020027);
`MEM('o011046, 16'o000017);
`MEM('o011050, 16'o001420);
`MEM('o011052, 16'o020027);
`MEM('o011054, 16'o000020);
`MEM('o011056, 16'o001032);
`MEM('o011060, 16'o016700);
`MEM('o011062, 16'o013102);
`MEM('o011064, 16'o005200);
`MEM('o011066, 16'o010067);
`MEM('o011070, 16'o013074);
`MEM('o011072, 16'o004767);
`MEM('o011074, 16'o177442);
`MEM('o011076, 16'o010065);
`MEM('o011100, 16'o177774);
`MEM('o011102, 16'o066565);
`MEM('o011104, 16'o177774);
`MEM('o011106, 16'o177776);
`MEM('o011110, 16'o000420);
`MEM('o011112, 16'o016700);
`MEM('o011114, 16'o013050);
`MEM('o011116, 16'o005200);
`MEM('o011120, 16'o010067);
`MEM('o011122, 16'o013042);
`MEM('o011124, 16'o004767);
`MEM('o011126, 16'o177410);
`MEM('o011130, 16'o010065);
`MEM('o011132, 16'o177774);
`MEM('o011134, 16'o166565);
`MEM('o011136, 16'o177774);
`MEM('o011140, 16'o177776);
`MEM('o011142, 16'o000403);
`MEM('o011144, 16'o016500);
`MEM('o011146, 16'o177776);
`MEM('o011150, 16'o000401);
`MEM('o011152, 16'o000727);
`MEM('o011154, 16'o010506);
`MEM('o011156, 16'o012605);
`MEM('o011160, 16'o000207);
`MEM('o011162, 16'o010546);
`MEM('o011164, 16'o010605);
`MEM('o011166, 16'o062706);
`MEM('o011170, 16'o177774);
`MEM('o011172, 16'o004767);
`MEM('o011174, 16'o177576);
`MEM('o011176, 16'o010065);
`MEM('o011200, 16'o177776);
`MEM('o011202, 16'o116700);
`MEM('o011204, 16'o007442);
`MEM('o011206, 16'o105700);
`MEM('o011210, 16'o001404);
`MEM('o011212, 16'o012700);
`MEM('o011214, 16'o177777);
`MEM('o011216, 16'o000167);
`MEM('o011220, 16'o000462);
`MEM('o011222, 16'o016700);
`MEM('o011224, 16'o012740);
`MEM('o011226, 16'o111000);
`MEM('o011230, 16'o042700);
`MEM('o011232, 16'o177400);
`MEM('o011234, 16'o062700);
`MEM('o011236, 16'o177753);
`MEM('o011240, 16'o020027);
`MEM('o011242, 16'o000005);
`MEM('o011244, 16'o101402);
`MEM('o011246, 16'o000167);
`MEM('o011250, 16'o000420);
`MEM('o011252, 16'o006300);
`MEM('o011254, 16'o062700);
`MEM('o011256, 16'o024320);
`MEM('o011260, 16'o011000);
`MEM('o011262, 16'o000110);
`MEM('o011264, 16'o016700);
`MEM('o011266, 16'o012676);
`MEM('o011270, 16'o005200);
`MEM('o011272, 16'o010067);
`MEM('o011274, 16'o012670);
`MEM('o011276, 16'o004767);
`MEM('o011300, 16'o177472);
`MEM('o011302, 16'o010065);
`MEM('o011304, 16'o177774);
`MEM('o011306, 16'o112700);
`MEM('o011310, 16'o000001);
`MEM('o011312, 16'o026565);
`MEM('o011314, 16'o177776);
`MEM('o011316, 16'o177774);
`MEM('o011320, 16'o001401);
`MEM('o011322, 16'o105000);
`MEM('o011324, 16'o005001);
`MEM('o011326, 16'o150001);
`MEM('o011330, 16'o010165);
`MEM('o011332, 16'o177776);
`MEM('o011334, 16'o000561);
`MEM('o011336, 16'o016700);
`MEM('o011340, 16'o012624);
`MEM('o011342, 16'o005200);
`MEM('o011344, 16'o010067);
`MEM('o011346, 16'o012616);
`MEM('o011350, 16'o004767);
`MEM('o011352, 16'o177420);
`MEM('o011354, 16'o010065);
`MEM('o011356, 16'o177774);
`MEM('o011360, 16'o016500);
`MEM('o011362, 16'o177774);
`MEM('o011364, 16'o016501);
`MEM('o011366, 16'o177776);
`MEM('o011370, 16'o074100);
`MEM('o011372, 16'o010001);
`MEM('o011374, 16'o005401);
`MEM('o011376, 16'o050100);
`MEM('o011400, 16'o000241);
`MEM('o011402, 16'o006000);
`MEM('o011404, 16'o072027);
`MEM('o011406, 16'o177762);
`MEM('o011410, 16'o005001);
`MEM('o011412, 16'o150001);
`MEM('o011414, 16'o010165);
`MEM('o011416, 16'o177776);
`MEM('o011420, 16'o000527);
`MEM('o011422, 16'o016700);
`MEM('o011424, 16'o012540);
`MEM('o011426, 16'o005200);
`MEM('o011430, 16'o010067);
`MEM('o011432, 16'o012532);
`MEM('o011434, 16'o004767);
`MEM('o011436, 16'o177334);
`MEM('o011440, 16'o010065);
`MEM('o011442, 16'o177774);
`MEM('o011444, 16'o112700);
`MEM('o011446, 16'o000001);
`MEM('o011450, 16'o026565);
`MEM('o011452, 16'o177776);
`MEM('o011454, 16'o177774);
`MEM('o011456, 16'o002401);
`MEM('o011460, 16'o105000);
`MEM('o011462, 16'o005001);
`MEM('o011464, 16'o150001);
`MEM('o011466, 16'o010165);
`MEM('o011470, 16'o177776);
`MEM('o011472, 16'o000502);
`MEM('o011474, 16'o016700);
`MEM('o011476, 16'o012466);
`MEM('o011500, 16'o005200);
`MEM('o011502, 16'o010067);
`MEM('o011504, 16'o012460);
`MEM('o011506, 16'o004767);
`MEM('o011510, 16'o177262);
`MEM('o011512, 16'o010065);
`MEM('o011514, 16'o177774);
`MEM('o011516, 16'o112700);
`MEM('o011520, 16'o000001);
`MEM('o011522, 16'o026565);
`MEM('o011524, 16'o177776);
`MEM('o011526, 16'o177774);
`MEM('o011530, 16'o003401);
`MEM('o011532, 16'o105000);
`MEM('o011534, 16'o005001);
`MEM('o011536, 16'o150001);
`MEM('o011540, 16'o010165);
`MEM('o011542, 16'o177776);
`MEM('o011544, 16'o000455);
`MEM('o011546, 16'o016700);
`MEM('o011550, 16'o012414);
`MEM('o011552, 16'o005200);
`MEM('o011554, 16'o010067);
`MEM('o011556, 16'o012406);
`MEM('o011560, 16'o004767);
`MEM('o011562, 16'o177210);
`MEM('o011564, 16'o010065);
`MEM('o011566, 16'o177774);
`MEM('o011570, 16'o112700);
`MEM('o011572, 16'o000001);
`MEM('o011574, 16'o026565);
`MEM('o011576, 16'o177776);
`MEM('o011600, 16'o177774);
`MEM('o011602, 16'o003001);
`MEM('o011604, 16'o105000);
`MEM('o011606, 16'o005001);
`MEM('o011610, 16'o150001);
`MEM('o011612, 16'o010165);
`MEM('o011614, 16'o177776);
`MEM('o011616, 16'o000430);
`MEM('o011620, 16'o016700);
`MEM('o011622, 16'o012342);
`MEM('o011624, 16'o005200);
`MEM('o011626, 16'o010067);
`MEM('o011630, 16'o012334);
`MEM('o011632, 16'o004767);
`MEM('o011634, 16'o177136);
`MEM('o011636, 16'o010065);
`MEM('o011640, 16'o177774);
`MEM('o011642, 16'o112700);
`MEM('o011644, 16'o000001);
`MEM('o011646, 16'o026565);
`MEM('o011650, 16'o177776);
`MEM('o011652, 16'o177774);
`MEM('o011654, 16'o002001);
`MEM('o011656, 16'o105000);
`MEM('o011660, 16'o005001);
`MEM('o011662, 16'o150001);
`MEM('o011664, 16'o010165);
`MEM('o011666, 16'o177776);
`MEM('o011670, 16'o000403);
`MEM('o011672, 16'o016500);
`MEM('o011674, 16'o177776);
`MEM('o011676, 16'o000402);
`MEM('o011700, 16'o000167);
`MEM('o011702, 16'o177316);
`MEM('o011704, 16'o010506);
`MEM('o011706, 16'o012605);
`MEM('o011710, 16'o000207);
`MEM('o011712, 16'o010546);
`MEM('o011714, 16'o010605);
`MEM('o011716, 16'o062706);
`MEM('o011720, 16'o177772);
`MEM('o011722, 16'o005065);
`MEM('o011724, 16'o177776);
`MEM('o011726, 16'o000167);
`MEM('o011730, 16'o000360);
`MEM('o011732, 16'o016700);
`MEM('o011734, 16'o012230);
`MEM('o011736, 16'o111000);
`MEM('o011740, 16'o042700);
`MEM('o011742, 16'o177400);
`MEM('o011744, 16'o020027);
`MEM('o011746, 16'o000026);
`MEM('o011750, 16'o001450);
`MEM('o011752, 16'o020027);
`MEM('o011754, 16'o000044);
`MEM('o011756, 16'o001063);
`MEM('o011760, 16'o016700);
`MEM('o011762, 16'o012202);
`MEM('o011764, 16'o005200);
`MEM('o011766, 16'o010067);
`MEM('o011770, 16'o012174);
`MEM('o011772, 16'o016700);
`MEM('o011774, 16'o012170);
`MEM('o011776, 16'o010001);
`MEM('o012000, 16'o005201);
`MEM('o012002, 16'o010167);
`MEM('o012004, 16'o012160);
`MEM('o012006, 16'o111065);
`MEM('o012010, 16'o177775);
`MEM('o012012, 16'o000416);
`MEM('o012014, 16'o016700);
`MEM('o012016, 16'o012146);
`MEM('o012020, 16'o010001);
`MEM('o012022, 16'o005201);
`MEM('o012024, 16'o010167);
`MEM('o012026, 16'o012136);
`MEM('o012030, 16'o111000);
`MEM('o012032, 16'o042700);
`MEM('o012034, 16'o177400);
`MEM('o012036, 16'o010046);
`MEM('o012040, 16'o004767);
`MEM('o012042, 16'o166744);
`MEM('o012044, 16'o062706);
`MEM('o012046, 16'o000002);
`MEM('o012050, 16'o116500);
`MEM('o012052, 16'o177775);
`MEM('o012054, 16'o110001);
`MEM('o012056, 16'o105301);
`MEM('o012060, 16'o110165);
`MEM('o012062, 16'o177775);
`MEM('o012064, 16'o105700);
`MEM('o012066, 16'o001352);
`MEM('o012070, 16'o000440);
`MEM('o012072, 16'o016700);
`MEM('o012074, 16'o012070);
`MEM('o012076, 16'o005200);
`MEM('o012100, 16'o010067);
`MEM('o012102, 16'o012062);
`MEM('o012104, 16'o004767);
`MEM('o012106, 16'o177052);
`MEM('o012110, 16'o010065);
`MEM('o012112, 16'o177776);
`MEM('o012114, 16'o116700);
`MEM('o012116, 16'o006530);
`MEM('o012120, 16'o105700);
`MEM('o012122, 16'o001422);
`MEM('o012124, 16'o000516);
`MEM('o012126, 16'o004767);
`MEM('o012130, 16'o177030);
`MEM('o012132, 16'o010065);
`MEM('o012134, 16'o177772);
`MEM('o012136, 16'o116700);
`MEM('o012140, 16'o006506);
`MEM('o012142, 16'o105700);
`MEM('o012144, 16'o001103);
`MEM('o012146, 16'o016546);
`MEM('o012150, 16'o177776);
`MEM('o012152, 16'o016546);
`MEM('o012154, 16'o177772);
`MEM('o012156, 16'o004767);
`MEM('o012160, 16'o170052);
`MEM('o012162, 16'o062706);
`MEM('o012164, 16'o000004);
`MEM('o012166, 16'o000401);
`MEM('o012170, 16'o000240);
`MEM('o012172, 16'o016700);
`MEM('o012174, 16'o011770);
`MEM('o012176, 16'o111000);
`MEM('o012200, 16'o120027);
`MEM('o012202, 16'o000015);
`MEM('o012204, 16'o001022);
`MEM('o012206, 16'o016700);
`MEM('o012210, 16'o011754);
`MEM('o012212, 16'o005200);
`MEM('o012214, 16'o010067);
`MEM('o012216, 16'o011746);
`MEM('o012220, 16'o016700);
`MEM('o012222, 16'o011742);
`MEM('o012224, 16'o111000);
`MEM('o012226, 16'o120027);
`MEM('o012230, 16'o000016);
`MEM('o012232, 16'o001452);
`MEM('o012234, 16'o016700);
`MEM('o012236, 16'o011726);
`MEM('o012240, 16'o111000);
`MEM('o012242, 16'o120027);
`MEM('o012244, 16'o000045);
`MEM('o012246, 16'o001021);
`MEM('o012250, 16'o000443);
`MEM('o012252, 16'o016700);
`MEM('o012254, 16'o011710);
`MEM('o012256, 16'o111000);
`MEM('o012260, 16'o120027);
`MEM('o012262, 16'o000016);
`MEM('o012264, 16'o001412);
`MEM('o012266, 16'o016700);
`MEM('o012270, 16'o011674);
`MEM('o012272, 16'o111000);
`MEM('o012274, 16'o120027);
`MEM('o012276, 16'o000045);
`MEM('o012300, 16'o001404);
`MEM('o012302, 16'o112767);
`MEM('o012304, 16'o000024);
`MEM('o012306, 16'o006340);
`MEM('o012310, 16'o000424);
`MEM('o012312, 16'o016700);
`MEM('o012314, 16'o011650);
`MEM('o012316, 16'o111000);
`MEM('o012320, 16'o120027);
`MEM('o012322, 16'o000016);
`MEM('o012324, 16'o001410);
`MEM('o012326, 16'o016700);
`MEM('o012330, 16'o011634);
`MEM('o012332, 16'o111000);
`MEM('o012334, 16'o120027);
`MEM('o012336, 16'o000045);
`MEM('o012340, 16'o001402);
`MEM('o012342, 16'o000167);
`MEM('o012344, 16'o177364);
`MEM('o012346, 16'o004767);
`MEM('o012350, 16'o166566);
`MEM('o012352, 16'o000403);
`MEM('o012354, 16'o000240);
`MEM('o012356, 16'o000401);
`MEM('o012360, 16'o000240);
`MEM('o012362, 16'o010506);
`MEM('o012364, 16'o012605);
`MEM('o012366, 16'o000207);
`MEM('o012370, 16'o010546);
`MEM('o012372, 16'o010605);
`MEM('o012374, 16'o062706);
`MEM('o012376, 16'o177772);
`MEM('o012400, 16'o112765);
`MEM('o012402, 16'o000001);
`MEM('o012404, 16'o177776);
`MEM('o012406, 16'o016700);
`MEM('o012410, 16'o011554);
`MEM('o012412, 16'o111000);
`MEM('o012414, 16'o120027);
`MEM('o012416, 16'o000044);
`MEM('o012420, 16'o001046);
`MEM('o012422, 16'o016700);
`MEM('o012424, 16'o011540);
`MEM('o012426, 16'o005200);
`MEM('o012430, 16'o010067);
`MEM('o012432, 16'o011532);
`MEM('o012434, 16'o016700);
`MEM('o012436, 16'o011526);
`MEM('o012440, 16'o010001);
`MEM('o012442, 16'o005201);
`MEM('o012444, 16'o010167);
`MEM('o012446, 16'o011516);
`MEM('o012450, 16'o111065);
`MEM('o012452, 16'o177777);
`MEM('o012454, 16'o000416);
`MEM('o012456, 16'o016700);
`MEM('o012460, 16'o011504);
`MEM('o012462, 16'o010001);
`MEM('o012464, 16'o005201);
`MEM('o012466, 16'o010167);
`MEM('o012470, 16'o011474);
`MEM('o012472, 16'o111000);
`MEM('o012474, 16'o042700);
`MEM('o012476, 16'o177400);
`MEM('o012500, 16'o010046);
`MEM('o012502, 16'o004767);
`MEM('o012504, 16'o166302);
`MEM('o012506, 16'o062706);
`MEM('o012510, 16'o000002);
`MEM('o012512, 16'o116500);
`MEM('o012514, 16'o177777);
`MEM('o012516, 16'o110001);
`MEM('o012520, 16'o105301);
`MEM('o012522, 16'o110165);
`MEM('o012524, 16'o177777);
`MEM('o012526, 16'o105700);
`MEM('o012530, 16'o001352);
`MEM('o012532, 16'o105065);
`MEM('o012534, 16'o177776);
`MEM('o012536, 16'o016700);
`MEM('o012540, 16'o011424);
`MEM('o012542, 16'o111000);
`MEM('o012544, 16'o042700);
`MEM('o012546, 16'o177400);
`MEM('o012550, 16'o020027);
`MEM('o012552, 16'o000033);
`MEM('o012554, 16'o001466);
`MEM('o012556, 16'o020027);
`MEM('o012560, 16'o000043);
`MEM('o012562, 16'o001156);
`MEM('o012564, 16'o016700);
`MEM('o012566, 16'o011376);
`MEM('o012570, 16'o005200);
`MEM('o012572, 16'o010067);
`MEM('o012574, 16'o011370);
`MEM('o012576, 16'o105765);
`MEM('o012600, 16'o177776);
`MEM('o012602, 16'o001422);
`MEM('o012604, 16'o016700);
`MEM('o012606, 16'o011356);
`MEM('o012610, 16'o111000);
`MEM('o012612, 16'o042700);
`MEM('o012614, 16'o177400);
`MEM('o012616, 16'o062700);
`MEM('o012620, 16'o000101);
`MEM('o012622, 16'o010046);
`MEM('o012624, 16'o004767);
`MEM('o012626, 16'o166160);
`MEM('o012630, 16'o062706);
`MEM('o012632, 16'o000002);
`MEM('o012634, 16'o012746);
`MEM('o012636, 16'o000072);
`MEM('o012640, 16'o004767);
`MEM('o012642, 16'o166144);
`MEM('o012644, 16'o062706);
`MEM('o012646, 16'o000002);
`MEM('o012650, 16'o004767);
`MEM('o012652, 16'o167654);
`MEM('o012654, 16'o010065);
`MEM('o012656, 16'o177774);
`MEM('o012660, 16'o116700);
`MEM('o012662, 16'o005764);
`MEM('o012664, 16'o105700);
`MEM('o012666, 16'o001402);
`MEM('o012670, 16'o000167);
`MEM('o012672, 16'o000330);
`MEM('o012674, 16'o016700);
`MEM('o012676, 16'o011266);
`MEM('o012700, 16'o010001);
`MEM('o012702, 16'o005201);
`MEM('o012704, 16'o010167);
`MEM('o012706, 16'o011256);
`MEM('o012710, 16'o111000);
`MEM('o012712, 16'o042700);
`MEM('o012714, 16'o177400);
`MEM('o012716, 16'o006300);
`MEM('o012720, 16'o062700);
`MEM('o012722, 16'o022000);
`MEM('o012724, 16'o016510);
`MEM('o012726, 16'o177774);
`MEM('o012730, 16'o000477);
`MEM('o012732, 16'o016700);
`MEM('o012734, 16'o011230);
`MEM('o012736, 16'o005200);
`MEM('o012740, 16'o010067);
`MEM('o012742, 16'o011222);
`MEM('o012744, 16'o004767);
`MEM('o012746, 16'o174610);
`MEM('o012750, 16'o010065);
`MEM('o012752, 16'o177772);
`MEM('o012754, 16'o116700);
`MEM('o012756, 16'o005670);
`MEM('o012760, 16'o105700);
`MEM('o012762, 16'o001122);
`MEM('o012764, 16'o026527);
`MEM('o012766, 16'o177772);
`MEM('o012770, 16'o000037);
`MEM('o012772, 16'o003404);
`MEM('o012774, 16'o112767);
`MEM('o012776, 16'o000003);
`MEM('o013000, 16'o005646);
`MEM('o013002, 16'o000517);
`MEM('o013004, 16'o105765);
`MEM('o013006, 16'o177776);
`MEM('o013010, 16'o001423);
`MEM('o013012, 16'o012746);
`MEM('o013014, 16'o024334);
`MEM('o013016, 16'o004767);
`MEM('o013020, 16'o166542);
`MEM('o013022, 16'o062706);
`MEM('o013024, 16'o000002);
`MEM('o013026, 16'o005046);
`MEM('o013030, 16'o016546);
`MEM('o013032, 16'o177772);
`MEM('o013034, 16'o004767);
`MEM('o013036, 16'o167174);
`MEM('o013040, 16'o062706);
`MEM('o013042, 16'o000004);
`MEM('o013044, 16'o012746);
`MEM('o013046, 16'o024337);
`MEM('o013050, 16'o004767);
`MEM('o013052, 16'o166510);
`MEM('o013054, 16'o062706);
`MEM('o013056, 16'o000002);
`MEM('o013060, 16'o004767);
`MEM('o013062, 16'o167444);
`MEM('o013064, 16'o010065);
`MEM('o013066, 16'o177774);
`MEM('o013070, 16'o116700);
`MEM('o013072, 16'o005554);
`MEM('o013074, 16'o105700);
`MEM('o013076, 16'o001056);
`MEM('o013100, 16'o016500);
`MEM('o013102, 16'o177772);
`MEM('o013104, 16'o006300);
`MEM('o013106, 16'o062700);
`MEM('o013110, 16'o022064);
`MEM('o013112, 16'o016510);
`MEM('o013114, 16'o177774);
`MEM('o013116, 16'o000404);
`MEM('o013120, 16'o112767);
`MEM('o013122, 16'o000024);
`MEM('o013124, 16'o005522);
`MEM('o013126, 16'o000445);
`MEM('o013130, 16'o016700);
`MEM('o013132, 16'o011032);
`MEM('o013134, 16'o111000);
`MEM('o013136, 16'o042700);
`MEM('o013140, 16'o177400);
`MEM('o013142, 16'o020027);
`MEM('o013144, 16'o000045);
`MEM('o013146, 16'o001434);
`MEM('o013150, 16'o020027);
`MEM('o013152, 16'o000045);
`MEM('o013154, 16'o003015);
`MEM('o013156, 16'o020027);
`MEM('o013160, 16'o000015);
`MEM('o013162, 16'o001404);
`MEM('o013164, 16'o020027);
`MEM('o013166, 16'o000016);
`MEM('o013170, 16'o001423);
`MEM('o013172, 16'o000406);
`MEM('o013174, 16'o016700);
`MEM('o013176, 16'o010766);
`MEM('o013200, 16'o005200);
`MEM('o013202, 16'o010067);
`MEM('o013204, 16'o010760);
`MEM('o013206, 16'o000404);
`MEM('o013210, 16'o112767);
`MEM('o013212, 16'o000024);
`MEM('o013214, 16'o005432);
`MEM('o013216, 16'o000411);
`MEM('o013220, 16'o000167);
`MEM('o013222, 16'o177154);
`MEM('o013224, 16'o000240);
`MEM('o013226, 16'o000405);
`MEM('o013230, 16'o000240);
`MEM('o013232, 16'o000403);
`MEM('o013234, 16'o000240);
`MEM('o013236, 16'o000401);
`MEM('o013240, 16'o000240);
`MEM('o013242, 16'o010506);
`MEM('o013244, 16'o012605);
`MEM('o013246, 16'o000207);
`MEM('o013250, 16'o010546);
`MEM('o013252, 16'o010605);
`MEM('o013254, 16'o062706);
`MEM('o013256, 16'o177774);
`MEM('o013260, 16'o016700);
`MEM('o013262, 16'o010702);
`MEM('o013264, 16'o010001);
`MEM('o013266, 16'o005201);
`MEM('o013270, 16'o010167);
`MEM('o013272, 16'o010672);
`MEM('o013274, 16'o111000);
`MEM('o013276, 16'o005001);
`MEM('o013300, 16'o150001);
`MEM('o013302, 16'o010165);
`MEM('o013304, 16'o177776);
`MEM('o013306, 16'o016700);
`MEM('o013310, 16'o010654);
`MEM('o013312, 16'o111000);
`MEM('o013314, 16'o120027);
`MEM('o013316, 16'o000030);
`MEM('o013320, 16'o001404);
`MEM('o013322, 16'o112767);
`MEM('o013324, 16'o000022);
`MEM('o013326, 16'o005320);
`MEM('o013330, 16'o000426);
`MEM('o013332, 16'o016700);
`MEM('o013334, 16'o010630);
`MEM('o013336, 16'o005200);
`MEM('o013340, 16'o010067);
`MEM('o013342, 16'o010622);
`MEM('o013344, 16'o004767);
`MEM('o013346, 16'o175612);
`MEM('o013350, 16'o010065);
`MEM('o013352, 16'o177774);
`MEM('o013354, 16'o116700);
`MEM('o013356, 16'o005270);
`MEM('o013360, 16'o105700);
`MEM('o013362, 16'o001010);
`MEM('o013364, 16'o016500);
`MEM('o013366, 16'o177776);
`MEM('o013370, 16'o006300);
`MEM('o013372, 16'o062700);
`MEM('o013374, 16'o022000);
`MEM('o013376, 16'o016510);
`MEM('o013400, 16'o177774);
`MEM('o013402, 16'o000401);
`MEM('o013404, 16'o000240);
`MEM('o013406, 16'o010506);
`MEM('o013410, 16'o012605);
`MEM('o013412, 16'o000207);
`MEM('o013414, 16'o010546);
`MEM('o013416, 16'o010605);
`MEM('o013420, 16'o062706);
`MEM('o013422, 16'o177774);
`MEM('o013424, 16'o004767);
`MEM('o013426, 16'o174130);
`MEM('o013430, 16'o010065);
`MEM('o013432, 16'o177776);
`MEM('o013434, 16'o116700);
`MEM('o013436, 16'o005210);
`MEM('o013440, 16'o105700);
`MEM('o013442, 16'o001047);
`MEM('o013444, 16'o026527);
`MEM('o013446, 16'o177776);
`MEM('o013450, 16'o000037);
`MEM('o013452, 16'o003404);
`MEM('o013454, 16'o112767);
`MEM('o013456, 16'o000003);
`MEM('o013460, 16'o005166);
`MEM('o013462, 16'o000442);
`MEM('o013464, 16'o016700);
`MEM('o013466, 16'o010476);
`MEM('o013470, 16'o111000);
`MEM('o013472, 16'o120027);
`MEM('o013474, 16'o000030);
`MEM('o013476, 16'o001404);
`MEM('o013500, 16'o112767);
`MEM('o013502, 16'o000022);
`MEM('o013504, 16'o005142);
`MEM('o013506, 16'o000430);
`MEM('o013510, 16'o016700);
`MEM('o013512, 16'o010452);
`MEM('o013514, 16'o005200);
`MEM('o013516, 16'o010067);
`MEM('o013520, 16'o010444);
`MEM('o013522, 16'o004767);
`MEM('o013524, 16'o175434);
`MEM('o013526, 16'o010065);
`MEM('o013530, 16'o177774);
`MEM('o013532, 16'o116700);
`MEM('o013534, 16'o005112);
`MEM('o013536, 16'o105700);
`MEM('o013540, 16'o001012);
`MEM('o013542, 16'o016500);
`MEM('o013544, 16'o177776);
`MEM('o013546, 16'o006300);
`MEM('o013550, 16'o062700);
`MEM('o013552, 16'o022064);
`MEM('o013554, 16'o016510);
`MEM('o013556, 16'o177774);
`MEM('o013560, 16'o000403);
`MEM('o013562, 16'o000240);
`MEM('o013564, 16'o000401);
`MEM('o013566, 16'o000240);
`MEM('o013570, 16'o010506);
`MEM('o013572, 16'o012605);
`MEM('o013574, 16'o000207);
`MEM('o013576, 16'o010546);
`MEM('o013600, 16'o010605);
`MEM('o013602, 16'o016700);
`MEM('o013604, 16'o010360);
`MEM('o013606, 16'o111000);
`MEM('o013610, 16'o042700);
`MEM('o013612, 16'o177400);
`MEM('o013614, 16'o020027);
`MEM('o013616, 16'o000033);
`MEM('o013620, 16'o001413);
`MEM('o013622, 16'o020027);
`MEM('o013624, 16'o000043);
`MEM('o013626, 16'o001020);
`MEM('o013630, 16'o016700);
`MEM('o013632, 16'o010332);
`MEM('o013634, 16'o005200);
`MEM('o013636, 16'o010067);
`MEM('o013640, 16'o010324);
`MEM('o013642, 16'o004767);
`MEM('o013644, 16'o177402);
`MEM('o013646, 16'o000414);
`MEM('o013650, 16'o016700);
`MEM('o013652, 16'o010312);
`MEM('o013654, 16'o005200);
`MEM('o013656, 16'o010067);
`MEM('o013660, 16'o010304);
`MEM('o013662, 16'o004767);
`MEM('o013664, 16'o177526);
`MEM('o013666, 16'o000404);
`MEM('o013670, 16'o112767);
`MEM('o013672, 16'o000016);
`MEM('o013674, 16'o004752);
`MEM('o013676, 16'o000240);
`MEM('o013700, 16'o000240);
`MEM('o013702, 16'o012605);
`MEM('o013704, 16'o000207);
`MEM('o013706, 16'o010546);
`MEM('o013710, 16'o010605);
`MEM('o013712, 16'o062706);
`MEM('o013714, 16'o177764);
`MEM('o013716, 16'o000167);
`MEM('o013720, 16'o002452);
`MEM('o013722, 16'o004767);
`MEM('o013724, 16'o165160);
`MEM('o013726, 16'o005700);
`MEM('o013730, 16'o001412);
`MEM('o013732, 16'o004767);
`MEM('o013734, 16'o165112);
`MEM('o013736, 16'o020027);
`MEM('o013740, 16'o000033);
`MEM('o013742, 16'o001005);
`MEM('o013744, 16'o112767);
`MEM('o013746, 16'o000026);
`MEM('o013750, 16'o004676);
`MEM('o013752, 16'o000167);
`MEM('o013754, 16'o002436);
`MEM('o013756, 16'o016700);
`MEM('o013760, 16'o010204);
`MEM('o013762, 16'o111000);
`MEM('o013764, 16'o042700);
`MEM('o013766, 16'o177400);
`MEM('o013770, 16'o020027);
`MEM('o013772, 16'o000043);
`MEM('o013774, 16'o101402);
`MEM('o013776, 16'o000167);
`MEM('o014000, 16'o002330);
`MEM('o014002, 16'o006300);
`MEM('o014004, 16'o062700);
`MEM('o014006, 16'o024342);
`MEM('o014010, 16'o011000);
`MEM('o014012, 16'o000110);
`MEM('o014014, 16'o016700);
`MEM('o014016, 16'o010146);
`MEM('o014020, 16'o005200);
`MEM('o014022, 16'o010067);
`MEM('o014024, 16'o010140);
`MEM('o014026, 16'o004767);
`MEM('o014030, 16'o175130);
`MEM('o014032, 16'o010065);
`MEM('o014034, 16'o177766);
`MEM('o014036, 16'o116700);
`MEM('o014040, 16'o004606);
`MEM('o014042, 16'o105700);
`MEM('o014044, 16'o001402);
`MEM('o014046, 16'o000167);
`MEM('o014050, 16'o002270);
`MEM('o014052, 16'o016546);
`MEM('o014054, 16'o177766);
`MEM('o014056, 16'o004767);
`MEM('o014060, 16'o171470);
`MEM('o014062, 16'o062706);
`MEM('o014064, 16'o000002);
`MEM('o014066, 16'o010065);
`MEM('o014070, 16'o177764);
`MEM('o014072, 16'o016546);
`MEM('o014074, 16'o177764);
`MEM('o014076, 16'o004767);
`MEM('o014100, 16'o171362);
`MEM('o014102, 16'o062706);
`MEM('o014104, 16'o000002);
`MEM('o014106, 16'o026500);
`MEM('o014110, 16'o177766);
`MEM('o014112, 16'o001405);
`MEM('o014114, 16'o112767);
`MEM('o014116, 16'o000020);
`MEM('o014120, 16'o004526);
`MEM('o014122, 16'o000167);
`MEM('o014124, 16'o002232);
`MEM('o014126, 16'o016567);
`MEM('o014130, 16'o177764);
`MEM('o014132, 16'o010030);
`MEM('o014134, 16'o016700);
`MEM('o014136, 16'o010024);
`MEM('o014140, 16'o062700);
`MEM('o014142, 16'o000003);
`MEM('o014144, 16'o010067);
`MEM('o014146, 16'o010016);
`MEM('o014150, 16'o000167);
`MEM('o014152, 16'o002204);
`MEM('o014154, 16'o016700);
`MEM('o014156, 16'o010006);
`MEM('o014160, 16'o005200);
`MEM('o014162, 16'o010067);
`MEM('o014164, 16'o010000);
`MEM('o014166, 16'o004767);
`MEM('o014170, 16'o174770);
`MEM('o014172, 16'o010065);
`MEM('o014174, 16'o177766);
`MEM('o014176, 16'o116700);
`MEM('o014200, 16'o004446);
`MEM('o014202, 16'o105700);
`MEM('o014204, 16'o001402);
`MEM('o014206, 16'o000167);
`MEM('o014210, 16'o002134);
`MEM('o014212, 16'o016546);
`MEM('o014214, 16'o177766);
`MEM('o014216, 16'o004767);
`MEM('o014220, 16'o171330);
`MEM('o014222, 16'o062706);
`MEM('o014224, 16'o000002);
`MEM('o014226, 16'o010065);
`MEM('o014230, 16'o177764);
`MEM('o014232, 16'o016546);
`MEM('o014234, 16'o177764);
`MEM('o014236, 16'o004767);
`MEM('o014240, 16'o171222);
`MEM('o014242, 16'o062706);
`MEM('o014244, 16'o000002);
`MEM('o014246, 16'o026500);
`MEM('o014250, 16'o177766);
`MEM('o014252, 16'o001405);
`MEM('o014254, 16'o112767);
`MEM('o014256, 16'o000020);
`MEM('o014260, 16'o004366);
`MEM('o014262, 16'o000167);
`MEM('o014264, 16'o002072);
`MEM('o014266, 16'o116700);
`MEM('o014270, 16'o007712);
`MEM('o014272, 16'o120027);
`MEM('o014274, 16'o000003);
`MEM('o014276, 16'o101405);
`MEM('o014300, 16'o112767);
`MEM('o014302, 16'o000006);
`MEM('o014304, 16'o004342);
`MEM('o014306, 16'o000167);
`MEM('o014310, 16'o002046);
`MEM('o014312, 16'o116700);
`MEM('o014314, 16'o007666);
`MEM('o014316, 16'o110001);
`MEM('o014320, 16'o105201);
`MEM('o014322, 16'o110167);
`MEM('o014324, 16'o007656);
`MEM('o014326, 16'o042700);
`MEM('o014330, 16'o177400);
`MEM('o014332, 16'o016701);
`MEM('o014334, 16'o007626);
`MEM('o014336, 16'o006300);
`MEM('o014340, 16'o062700);
`MEM('o014342, 16'o024170);
`MEM('o014344, 16'o010110);
`MEM('o014346, 16'o116700);
`MEM('o014350, 16'o007632);
`MEM('o014352, 16'o110001);
`MEM('o014354, 16'o105201);
`MEM('o014356, 16'o110167);
`MEM('o014360, 16'o007622);
`MEM('o014362, 16'o042700);
`MEM('o014364, 16'o177400);
`MEM('o014366, 16'o016701);
`MEM('o014370, 16'o007574);
`MEM('o014372, 16'o006300);
`MEM('o014374, 16'o062700);
`MEM('o014376, 16'o024170);
`MEM('o014400, 16'o010110);
`MEM('o014402, 16'o016567);
`MEM('o014404, 16'o177764);
`MEM('o014406, 16'o007554);
`MEM('o014410, 16'o016700);
`MEM('o014412, 16'o007550);
`MEM('o014414, 16'o062700);
`MEM('o014416, 16'o000003);
`MEM('o014420, 16'o010067);
`MEM('o014422, 16'o007542);
`MEM('o014424, 16'o000167);
`MEM('o014426, 16'o001730);
`MEM('o014430, 16'o116700);
`MEM('o014432, 16'o007550);
`MEM('o014434, 16'o120027);
`MEM('o014436, 16'o000001);
`MEM('o014440, 16'o101005);
`MEM('o014442, 16'o112767);
`MEM('o014444, 16'o000007);
`MEM('o014446, 16'o004200);
`MEM('o014450, 16'o000167);
`MEM('o014452, 16'o001704);
`MEM('o014454, 16'o116700);
`MEM('o014456, 16'o007524);
`MEM('o014460, 16'o105300);
`MEM('o014462, 16'o110067);
`MEM('o014464, 16'o007516);
`MEM('o014466, 16'o116700);
`MEM('o014470, 16'o007512);
`MEM('o014472, 16'o042700);
`MEM('o014474, 16'o177400);
`MEM('o014476, 16'o006300);
`MEM('o014500, 16'o062700);
`MEM('o014502, 16'o024170);
`MEM('o014504, 16'o011000);
`MEM('o014506, 16'o010067);
`MEM('o014510, 16'o007454);
`MEM('o014512, 16'o116700);
`MEM('o014514, 16'o007466);
`MEM('o014516, 16'o105300);
`MEM('o014520, 16'o110067);
`MEM('o014522, 16'o007460);
`MEM('o014524, 16'o116700);
`MEM('o014526, 16'o007454);
`MEM('o014530, 16'o042700);
`MEM('o014532, 16'o177400);
`MEM('o014534, 16'o006300);
`MEM('o014536, 16'o062700);
`MEM('o014540, 16'o024170);
`MEM('o014542, 16'o011000);
`MEM('o014544, 16'o010067);
`MEM('o014546, 16'o007414);
`MEM('o014550, 16'o000167);
`MEM('o014552, 16'o001604);
`MEM('o014554, 16'o016700);
`MEM('o014556, 16'o007406);
`MEM('o014560, 16'o005200);
`MEM('o014562, 16'o010067);
`MEM('o014564, 16'o007400);
`MEM('o014566, 16'o016700);
`MEM('o014570, 16'o007374);
`MEM('o014572, 16'o010001);
`MEM('o014574, 16'o005201);
`MEM('o014576, 16'o010167);
`MEM('o014600, 16'o007364);
`MEM('o014602, 16'o111000);
`MEM('o014604, 16'o120027);
`MEM('o014606, 16'o000043);
`MEM('o014610, 16'o001405);
`MEM('o014612, 16'o112767);
`MEM('o014614, 16'o000014);
`MEM('o014616, 16'o004030);
`MEM('o014620, 16'o000167);
`MEM('o014622, 16'o001534);
`MEM('o014624, 16'o016700);
`MEM('o014626, 16'o007336);
`MEM('o014630, 16'o111000);
`MEM('o014632, 16'o005001);
`MEM('o014634, 16'o150001);
`MEM('o014636, 16'o010165);
`MEM('o014640, 16'o177772);
`MEM('o014642, 16'o004767);
`MEM('o014644, 16'o176402);
`MEM('o014646, 16'o116700);
`MEM('o014650, 16'o003776);
`MEM('o014652, 16'o105700);
`MEM('o014654, 16'o001402);
`MEM('o014656, 16'o000167);
`MEM('o014660, 16'o001470);
`MEM('o014662, 16'o016700);
`MEM('o014664, 16'o007300);
`MEM('o014666, 16'o111000);
`MEM('o014670, 16'o120027);
`MEM('o014672, 16'o000004);
`MEM('o014674, 16'o001020);
`MEM('o014676, 16'o016700);
`MEM('o014700, 16'o007264);
`MEM('o014702, 16'o005200);
`MEM('o014704, 16'o010067);
`MEM('o014706, 16'o007256);
`MEM('o014710, 16'o004767);
`MEM('o014712, 16'o174246);
`MEM('o014714, 16'o010065);
`MEM('o014716, 16'o177770);
`MEM('o014720, 16'o016700);
`MEM('o014722, 16'o007242);
`MEM('o014724, 16'o111000);
`MEM('o014726, 16'o120027);
`MEM('o014730, 16'o000005);
`MEM('o014732, 16'o001020);
`MEM('o014734, 16'o000405);
`MEM('o014736, 16'o112767);
`MEM('o014740, 16'o000015);
`MEM('o014742, 16'o003704);
`MEM('o014744, 16'o000167);
`MEM('o014746, 16'o001410);
`MEM('o014750, 16'o016700);
`MEM('o014752, 16'o007212);
`MEM('o014754, 16'o005200);
`MEM('o014756, 16'o010067);
`MEM('o014760, 16'o007204);
`MEM('o014762, 16'o004767);
`MEM('o014764, 16'o174174);
`MEM('o014766, 16'o010065);
`MEM('o014770, 16'o177776);
`MEM('o014772, 16'o000403);
`MEM('o014774, 16'o012765);
`MEM('o014776, 16'o000001);
`MEM('o015000, 16'o177776);
`MEM('o015002, 16'o005765);
`MEM('o015004, 16'o177776);
`MEM('o015006, 16'o002007);
`MEM('o015010, 16'o012700);
`MEM('o015012, 16'o100001);
`MEM('o015014, 16'o166500);
`MEM('o015016, 16'o177776);
`MEM('o015020, 16'o026500);
`MEM('o015022, 16'o177770);
`MEM('o015024, 16'o002412);
`MEM('o015026, 16'o005765);
`MEM('o015030, 16'o177776);
`MEM('o015032, 16'o003414);
`MEM('o015034, 16'o012700);
`MEM('o015036, 16'o077777);
`MEM('o015040, 16'o166500);
`MEM('o015042, 16'o177776);
`MEM('o015044, 16'o026500);
`MEM('o015046, 16'o177770);
`MEM('o015050, 16'o003405);
`MEM('o015052, 16'o112767);
`MEM('o015054, 16'o000002);
`MEM('o015056, 16'o003570);
`MEM('o015060, 16'o000167);
`MEM('o015062, 16'o001274);
`MEM('o015064, 16'o116700);
`MEM('o015066, 16'o007154);
`MEM('o015070, 16'o120027);
`MEM('o015072, 16'o000011);
`MEM('o015074, 16'o101405);
`MEM('o015076, 16'o112767);
`MEM('o015100, 16'o000010);
`MEM('o015102, 16'o003544);
`MEM('o015104, 16'o000167);
`MEM('o015106, 16'o001250);
`MEM('o015110, 16'o116700);
`MEM('o015112, 16'o007130);
`MEM('o015114, 16'o110001);
`MEM('o015116, 16'o105201);
`MEM('o015120, 16'o110167);
`MEM('o015122, 16'o007120);
`MEM('o015124, 16'o042700);
`MEM('o015126, 16'o177400);
`MEM('o015130, 16'o016701);
`MEM('o015132, 16'o007030);
`MEM('o015134, 16'o006300);
`MEM('o015136, 16'o062700);
`MEM('o015140, 16'o024206);
`MEM('o015142, 16'o010110);
`MEM('o015144, 16'o116700);
`MEM('o015146, 16'o007074);
`MEM('o015150, 16'o110001);
`MEM('o015152, 16'o105201);
`MEM('o015154, 16'o110167);
`MEM('o015156, 16'o007064);
`MEM('o015160, 16'o042700);
`MEM('o015162, 16'o177400);
`MEM('o015164, 16'o016701);
`MEM('o015166, 16'o006776);
`MEM('o015170, 16'o006300);
`MEM('o015172, 16'o062700);
`MEM('o015174, 16'o024206);
`MEM('o015176, 16'o010110);
`MEM('o015200, 16'o116700);
`MEM('o015202, 16'o007040);
`MEM('o015204, 16'o110001);
`MEM('o015206, 16'o105201);
`MEM('o015210, 16'o110167);
`MEM('o015212, 16'o007030);
`MEM('o015214, 16'o042700);
`MEM('o015216, 16'o177400);
`MEM('o015220, 16'o016501);
`MEM('o015222, 16'o177770);
`MEM('o015224, 16'o006300);
`MEM('o015226, 16'o062700);
`MEM('o015230, 16'o024206);
`MEM('o015232, 16'o010110);
`MEM('o015234, 16'o116700);
`MEM('o015236, 16'o007004);
`MEM('o015240, 16'o110001);
`MEM('o015242, 16'o105201);
`MEM('o015244, 16'o110167);
`MEM('o015246, 16'o006774);
`MEM('o015250, 16'o042700);
`MEM('o015252, 16'o177400);
`MEM('o015254, 16'o016501);
`MEM('o015256, 16'o177776);
`MEM('o015260, 16'o006300);
`MEM('o015262, 16'o062700);
`MEM('o015264, 16'o024206);
`MEM('o015266, 16'o010110);
`MEM('o015270, 16'o116700);
`MEM('o015272, 16'o006750);
`MEM('o015274, 16'o110001);
`MEM('o015276, 16'o105201);
`MEM('o015300, 16'o110167);
`MEM('o015302, 16'o006740);
`MEM('o015304, 16'o042700);
`MEM('o015306, 16'o177400);
`MEM('o015310, 16'o016501);
`MEM('o015312, 16'o177772);
`MEM('o015314, 16'o006300);
`MEM('o015316, 16'o062700);
`MEM('o015320, 16'o024206);
`MEM('o015322, 16'o010110);
`MEM('o015324, 16'o000167);
`MEM('o015326, 16'o001030);
`MEM('o015330, 16'o016700);
`MEM('o015332, 16'o006632);
`MEM('o015334, 16'o005200);
`MEM('o015336, 16'o010067);
`MEM('o015340, 16'o006624);
`MEM('o015342, 16'o116700);
`MEM('o015344, 16'o006676);
`MEM('o015346, 16'o120027);
`MEM('o015350, 16'o000004);
`MEM('o015352, 16'o101005);
`MEM('o015354, 16'o112767);
`MEM('o015356, 16'o000011);
`MEM('o015360, 16'o003266);
`MEM('o015362, 16'o000167);
`MEM('o015364, 16'o000772);
`MEM('o015366, 16'o116700);
`MEM('o015370, 16'o006652);
`MEM('o015372, 16'o042700);
`MEM('o015374, 16'o177400);
`MEM('o015376, 16'o005300);
`MEM('o015400, 16'o006300);
`MEM('o015402, 16'o062700);
`MEM('o015404, 16'o024206);
`MEM('o015406, 16'o011000);
`MEM('o015410, 16'o010065);
`MEM('o015412, 16'o177772);
`MEM('o015414, 16'o016700);
`MEM('o015416, 16'o006546);
`MEM('o015420, 16'o010001);
`MEM('o015422, 16'o005201);
`MEM('o015424, 16'o010167);
`MEM('o015426, 16'o006536);
`MEM('o015430, 16'o111000);
`MEM('o015432, 16'o120027);
`MEM('o015434, 16'o000043);
`MEM('o015436, 16'o001405);
`MEM('o015440, 16'o112767);
`MEM('o015442, 16'o000012);
`MEM('o015444, 16'o003202);
`MEM('o015446, 16'o000167);
`MEM('o015450, 16'o000706);
`MEM('o015452, 16'o016700);
`MEM('o015454, 16'o006510);
`MEM('o015456, 16'o010001);
`MEM('o015460, 16'o005201);
`MEM('o015462, 16'o010167);
`MEM('o015464, 16'o006500);
`MEM('o015466, 16'o111000);
`MEM('o015470, 16'o042700);
`MEM('o015472, 16'o177400);
`MEM('o015474, 16'o026500);
`MEM('o015476, 16'o177772);
`MEM('o015500, 16'o001405);
`MEM('o015502, 16'o112767);
`MEM('o015504, 16'o000013);
`MEM('o015506, 16'o003140);
`MEM('o015510, 16'o000167);
`MEM('o015512, 16'o000644);
`MEM('o015514, 16'o116700);
`MEM('o015516, 16'o006524);
`MEM('o015520, 16'o042700);
`MEM('o015522, 16'o177400);
`MEM('o015524, 16'o062700);
`MEM('o015526, 16'o177776);
`MEM('o015530, 16'o006300);
`MEM('o015532, 16'o062700);
`MEM('o015534, 16'o024206);
`MEM('o015536, 16'o011000);
`MEM('o015540, 16'o010065);
`MEM('o015542, 16'o177776);
`MEM('o015544, 16'o016500);
`MEM('o015546, 16'o177772);
`MEM('o015550, 16'o006300);
`MEM('o015552, 16'o062700);
`MEM('o015554, 16'o022000);
`MEM('o015556, 16'o011000);
`MEM('o015560, 16'o016501);
`MEM('o015562, 16'o177776);
`MEM('o015564, 16'o060001);
`MEM('o015566, 16'o016500);
`MEM('o015570, 16'o177772);
`MEM('o015572, 16'o006300);
`MEM('o015574, 16'o062700);
`MEM('o015576, 16'o022000);
`MEM('o015600, 16'o010110);
`MEM('o015602, 16'o116700);
`MEM('o015604, 16'o006436);
`MEM('o015606, 16'o042700);
`MEM('o015610, 16'o177400);
`MEM('o015612, 16'o062700);
`MEM('o015614, 16'o177775);
`MEM('o015616, 16'o006300);
`MEM('o015620, 16'o062700);
`MEM('o015622, 16'o024206);
`MEM('o015624, 16'o011000);
`MEM('o015626, 16'o010065);
`MEM('o015630, 16'o177770);
`MEM('o015632, 16'o005765);
`MEM('o015634, 16'o177776);
`MEM('o015636, 16'o002011);
`MEM('o015640, 16'o016500);
`MEM('o015642, 16'o177772);
`MEM('o015644, 16'o006300);
`MEM('o015646, 16'o062700);
`MEM('o015650, 16'o022000);
`MEM('o015652, 16'o011000);
`MEM('o015654, 16'o026500);
`MEM('o015656, 16'o177770);
`MEM('o015660, 16'o003014);
`MEM('o015662, 16'o005765);
`MEM('o015664, 16'o177776);
`MEM('o015666, 16'o003421);
`MEM('o015670, 16'o016500);
`MEM('o015672, 16'o177772);
`MEM('o015674, 16'o006300);
`MEM('o015676, 16'o062700);
`MEM('o015700, 16'o022000);
`MEM('o015702, 16'o011000);
`MEM('o015704, 16'o026500);
`MEM('o015706, 16'o177770);
`MEM('o015710, 16'o002010);
`MEM('o015712, 16'o116700);
`MEM('o015714, 16'o006326);
`MEM('o015716, 16'o062700);
`MEM('o015720, 16'o177773);
`MEM('o015722, 16'o110067);
`MEM('o015724, 16'o006316);
`MEM('o015726, 16'o000167);
`MEM('o015730, 16'o000426);
`MEM('o015732, 16'o116700);
`MEM('o015734, 16'o006306);
`MEM('o015736, 16'o042700);
`MEM('o015740, 16'o177400);
`MEM('o015742, 16'o062700);
`MEM('o015744, 16'o177774);
`MEM('o015746, 16'o006300);
`MEM('o015750, 16'o062700);
`MEM('o015752, 16'o024206);
`MEM('o015754, 16'o011000);
`MEM('o015756, 16'o010067);
`MEM('o015760, 16'o006204);
`MEM('o015762, 16'o116700);
`MEM('o015764, 16'o006256);
`MEM('o015766, 16'o042700);
`MEM('o015770, 16'o177400);
`MEM('o015772, 16'o062700);
`MEM('o015774, 16'o177773);
`MEM('o015776, 16'o006300);
`MEM('o016000, 16'o062700);
`MEM('o016002, 16'o024206);
`MEM('o016004, 16'o011000);
`MEM('o016006, 16'o010067);
`MEM('o016010, 16'o006152);
`MEM('o016012, 16'o000167);
`MEM('o016014, 16'o000342);
`MEM('o016016, 16'o016700);
`MEM('o016020, 16'o006144);
`MEM('o016022, 16'o005200);
`MEM('o016024, 16'o010067);
`MEM('o016026, 16'o006136);
`MEM('o016030, 16'o004767);
`MEM('o016032, 16'o173126);
`MEM('o016034, 16'o010065);
`MEM('o016036, 16'o177774);
`MEM('o016040, 16'o116700);
`MEM('o016042, 16'o002604);
`MEM('o016044, 16'o105700);
`MEM('o016046, 16'o001404);
`MEM('o016050, 16'o112767);
`MEM('o016052, 16'o000017);
`MEM('o016054, 16'o002572);
`MEM('o016056, 16'o000540);
`MEM('o016060, 16'o005765);
`MEM('o016062, 16'o177774);
`MEM('o016064, 16'o001134);
`MEM('o016066, 16'o000405);
`MEM('o016070, 16'o016700);
`MEM('o016072, 16'o006072);
`MEM('o016074, 16'o005200);
`MEM('o016076, 16'o010067);
`MEM('o016100, 16'o006064);
`MEM('o016102, 16'o016700);
`MEM('o016104, 16'o006060);
`MEM('o016106, 16'o111000);
`MEM('o016110, 16'o120027);
`MEM('o016112, 16'o000045);
`MEM('o016114, 16'o001365);
`MEM('o016116, 16'o000520);
`MEM('o016120, 16'o016701);
`MEM('o016122, 16'o006040);
`MEM('o016124, 16'o016700);
`MEM('o016126, 16'o006034);
`MEM('o016130, 16'o111000);
`MEM('o016132, 16'o042700);
`MEM('o016134, 16'o177400);
`MEM('o016136, 16'o060100);
`MEM('o016140, 16'o010067);
`MEM('o016142, 16'o006020);
`MEM('o016144, 16'o016700);
`MEM('o016146, 16'o006014);
`MEM('o016150, 16'o111000);
`MEM('o016152, 16'o105700);
`MEM('o016154, 16'o001361);
`MEM('o016156, 16'o016700);
`MEM('o016160, 16'o006002);
`MEM('o016162, 16'o000524);
`MEM('o016164, 16'o016700);
`MEM('o016166, 16'o005776);
`MEM('o016170, 16'o005200);
`MEM('o016172, 16'o010067);
`MEM('o016174, 16'o005770);
`MEM('o016176, 16'o004767);
`MEM('o016200, 16'o175046);
`MEM('o016202, 16'o000466);
`MEM('o016204, 16'o016700);
`MEM('o016206, 16'o005756);
`MEM('o016210, 16'o005200);
`MEM('o016212, 16'o010067);
`MEM('o016214, 16'o005750);
`MEM('o016216, 16'o004767);
`MEM('o016220, 16'o175172);
`MEM('o016222, 16'o000456);
`MEM('o016224, 16'o016700);
`MEM('o016226, 16'o005736);
`MEM('o016230, 16'o005200);
`MEM('o016232, 16'o010067);
`MEM('o016234, 16'o005730);
`MEM('o016236, 16'o004767);
`MEM('o016240, 16'o175334);
`MEM('o016242, 16'o000446);
`MEM('o016244, 16'o016700);
`MEM('o016246, 16'o005716);
`MEM('o016250, 16'o005200);
`MEM('o016252, 16'o010067);
`MEM('o016254, 16'o005710);
`MEM('o016256, 16'o004767);
`MEM('o016260, 16'o173430);
`MEM('o016262, 16'o000436);
`MEM('o016264, 16'o016700);
`MEM('o016266, 16'o005676);
`MEM('o016270, 16'o005200);
`MEM('o016272, 16'o010067);
`MEM('o016274, 16'o005670);
`MEM('o016276, 16'o004767);
`MEM('o016300, 16'o174066);
`MEM('o016302, 16'o000426);
`MEM('o016304, 16'o112767);
`MEM('o016306, 16'o000023);
`MEM('o016310, 16'o002336);
`MEM('o016312, 16'o005000);
`MEM('o016314, 16'o000447);
`MEM('o016316, 16'o016700);
`MEM('o016320, 16'o005644);
`MEM('o016322, 16'o005200);
`MEM('o016324, 16'o010067);
`MEM('o016326, 16'o005636);
`MEM('o016330, 16'o000413);
`MEM('o016332, 16'o112767);
`MEM('o016334, 16'o000024);
`MEM('o016336, 16'o002310);
`MEM('o016340, 16'o000407);
`MEM('o016342, 16'o000240);
`MEM('o016344, 16'o000405);
`MEM('o016346, 16'o000240);
`MEM('o016350, 16'o000403);
`MEM('o016352, 16'o000240);
`MEM('o016354, 16'o000401);
`MEM('o016356, 16'o000240);
`MEM('o016360, 16'o116700);
`MEM('o016362, 16'o002264);
`MEM('o016364, 16'o105700);
`MEM('o016366, 16'o001402);
`MEM('o016370, 16'o005000);
`MEM('o016372, 16'o000420);
`MEM('o016374, 16'o016700);
`MEM('o016376, 16'o005566);
`MEM('o016400, 16'o111000);
`MEM('o016402, 16'o120027);
`MEM('o016404, 16'o000045);
`MEM('o016406, 16'o001402);
`MEM('o016410, 16'o000167);
`MEM('o016412, 16'o175306);
`MEM('o016414, 16'o016701);
`MEM('o016416, 16'o005544);
`MEM('o016420, 16'o016700);
`MEM('o016422, 16'o005540);
`MEM('o016424, 16'o111000);
`MEM('o016426, 16'o042700);
`MEM('o016430, 16'o177400);
`MEM('o016432, 16'o060100);
`MEM('o016434, 16'o010506);
`MEM('o016436, 16'o012605);
`MEM('o016440, 16'o000207);
`MEM('o016442, 16'o010546);
`MEM('o016444, 16'o010605);
`MEM('o016446, 16'o062706);
`MEM('o016450, 16'o177776);
`MEM('o016452, 16'o105067);
`MEM('o016454, 16'o005526);
`MEM('o016456, 16'o105067);
`MEM('o016460, 16'o005562);
`MEM('o016462, 16'o012767);
`MEM('o016464, 16'o022164);
`MEM('o016466, 16'o005474);
`MEM('o016470, 16'o000421);
`MEM('o016472, 16'o016700);
`MEM('o016474, 16'o005466);
`MEM('o016476, 16'o062700);
`MEM('o016500, 16'o000003);
`MEM('o016502, 16'o010067);
`MEM('o016504, 16'o005460);
`MEM('o016506, 16'o004767);
`MEM('o016510, 16'o175174);
`MEM('o016512, 16'o010065);
`MEM('o016514, 16'o177776);
`MEM('o016516, 16'o116700);
`MEM('o016520, 16'o002126);
`MEM('o016522, 16'o105700);
`MEM('o016524, 16'o001011);
`MEM('o016526, 16'o016567);
`MEM('o016530, 16'o177776);
`MEM('o016532, 16'o005430);
`MEM('o016534, 16'o016700);
`MEM('o016536, 16'o005424);
`MEM('o016540, 16'o111000);
`MEM('o016542, 16'o105700);
`MEM('o016544, 16'o001352);
`MEM('o016546, 16'o000401);
`MEM('o016550, 16'o000240);
`MEM('o016552, 16'o010506);
`MEM('o016554, 16'o012605);
`MEM('o016556, 16'o000207);
`MEM('o016560, 16'o010546);
`MEM('o016562, 16'o010605);
`MEM('o016564, 16'o062706);
`MEM('o016566, 16'o177776);
`MEM('o016570, 16'o016700);
`MEM('o016572, 16'o005372);
`MEM('o016574, 16'o111000);
`MEM('o016576, 16'o120027);
`MEM('o016600, 16'o000042);
`MEM('o016602, 16'o001012);
`MEM('o016604, 16'o016700);
`MEM('o016606, 16'o005356);
`MEM('o016610, 16'o010046);
`MEM('o016612, 16'o004767);
`MEM('o016614, 16'o166646);
`MEM('o016616, 16'o062706);
`MEM('o016620, 16'o000002);
`MEM('o016622, 16'o010065);
`MEM('o016624, 16'o177776);
`MEM('o016626, 16'o000402);
`MEM('o016630, 16'o005065);
`MEM('o016632, 16'o177776);
`MEM('o016634, 16'o012767);
`MEM('o016636, 16'o022164);
`MEM('o016640, 16'o005322);
`MEM('o016642, 16'o000412);
`MEM('o016644, 16'o016701);
`MEM('o016646, 16'o005314);
`MEM('o016650, 16'o016700);
`MEM('o016652, 16'o005310);
`MEM('o016654, 16'o111000);
`MEM('o016656, 16'o042700);
`MEM('o016660, 16'o177400);
`MEM('o016662, 16'o060100);
`MEM('o016664, 16'o010067);
`MEM('o016666, 16'o005274);
`MEM('o016670, 16'o016700);
`MEM('o016672, 16'o005270);
`MEM('o016674, 16'o111000);
`MEM('o016676, 16'o105700);
`MEM('o016700, 16'o001467);
`MEM('o016702, 16'o016700);
`MEM('o016704, 16'o005256);
`MEM('o016706, 16'o010046);
`MEM('o016710, 16'o004767);
`MEM('o016712, 16'o166550);
`MEM('o016714, 16'o062706);
`MEM('o016716, 16'o000002);
`MEM('o016720, 16'o026500);
`MEM('o016722, 16'o177776);
`MEM('o016724, 16'o003347);
`MEM('o016726, 16'o000454);
`MEM('o016730, 16'o016700);
`MEM('o016732, 16'o005230);
`MEM('o016734, 16'o010046);
`MEM('o016736, 16'o004767);
`MEM('o016740, 16'o166522);
`MEM('o016742, 16'o062706);
`MEM('o016744, 16'o000002);
`MEM('o016746, 16'o005046);
`MEM('o016750, 16'o010046);
`MEM('o016752, 16'o004767);
`MEM('o016754, 16'o163256);
`MEM('o016756, 16'o062706);
`MEM('o016760, 16'o000004);
`MEM('o016762, 16'o012746);
`MEM('o016764, 16'o000040);
`MEM('o016766, 16'o004767);
`MEM('o016770, 16'o162016);
`MEM('o016772, 16'o062706);
`MEM('o016774, 16'o000002);
`MEM('o016776, 16'o016700);
`MEM('o017000, 16'o005162);
`MEM('o017002, 16'o062700);
`MEM('o017004, 16'o000003);
`MEM('o017006, 16'o010046);
`MEM('o017010, 16'o004767);
`MEM('o017012, 16'o167442);
`MEM('o017014, 16'o062706);
`MEM('o017016, 16'o000002);
`MEM('o017020, 16'o116700);
`MEM('o017022, 16'o001624);
`MEM('o017024, 16'o105700);
`MEM('o017026, 16'o001022);
`MEM('o017030, 16'o004767);
`MEM('o017032, 16'o162104);
`MEM('o017034, 16'o016701);
`MEM('o017036, 16'o005124);
`MEM('o017040, 16'o016700);
`MEM('o017042, 16'o005120);
`MEM('o017044, 16'o111000);
`MEM('o017046, 16'o042700);
`MEM('o017050, 16'o177400);
`MEM('o017052, 16'o060100);
`MEM('o017054, 16'o010067);
`MEM('o017056, 16'o005104);
`MEM('o017060, 16'o016700);
`MEM('o017062, 16'o005100);
`MEM('o017064, 16'o111000);
`MEM('o017066, 16'o105700);
`MEM('o017070, 16'o001317);
`MEM('o017072, 16'o000401);
`MEM('o017074, 16'o000240);
`MEM('o017076, 16'o000240);
`MEM('o017100, 16'o010506);
`MEM('o017102, 16'o012605);
`MEM('o017104, 16'o000207);
`MEM('o017106, 16'o010546);
`MEM('o017110, 16'o010605);
`MEM('o017112, 16'o062706);
`MEM('o017114, 16'o177776);
`MEM('o017116, 16'o105065);
`MEM('o017120, 16'o177777);
`MEM('o017122, 16'o000415);
`MEM('o017124, 16'o005000);
`MEM('o017126, 16'o156500);
`MEM('o017130, 16'o177777);
`MEM('o017132, 16'o006300);
`MEM('o017134, 16'o062700);
`MEM('o017136, 16'o022000);
`MEM('o017140, 16'o005010);
`MEM('o017142, 16'o116500);
`MEM('o017144, 16'o177777);
`MEM('o017146, 16'o110001);
`MEM('o017150, 16'o105201);
`MEM('o017152, 16'o110165);
`MEM('o017154, 16'o177777);
`MEM('o017156, 16'o126527);
`MEM('o017160, 16'o177777);
`MEM('o017162, 16'o000031);
`MEM('o017164, 16'o101757);
`MEM('o017166, 16'o105065);
`MEM('o017170, 16'o177777);
`MEM('o017172, 16'o000415);
`MEM('o017174, 16'o005000);
`MEM('o017176, 16'o156500);
`MEM('o017200, 16'o177777);
`MEM('o017202, 16'o006300);
`MEM('o017204, 16'o062700);
`MEM('o017206, 16'o022064);
`MEM('o017210, 16'o005010);
`MEM('o017212, 16'o116500);
`MEM('o017214, 16'o177777);
`MEM('o017216, 16'o110001);
`MEM('o017220, 16'o105201);
`MEM('o017222, 16'o110165);
`MEM('o017224, 16'o177777);
`MEM('o017226, 16'o126527);
`MEM('o017230, 16'o177777);
`MEM('o017232, 16'o000037);
`MEM('o017234, 16'o101757);
`MEM('o017236, 16'o105067);
`MEM('o017240, 16'o004742);
`MEM('o017242, 16'o105067);
`MEM('o017244, 16'o004776);
`MEM('o017246, 16'o105067);
`MEM('o017250, 16'o002712);
`MEM('o017252, 16'o012767);
`MEM('o017254, 16'o022164);
`MEM('o017256, 16'o004704);
`MEM('o017260, 16'o000240);
`MEM('o017262, 16'o010506);
`MEM('o017264, 16'o012605);
`MEM('o017266, 16'o000207);
`MEM('o017270, 16'o010546);
`MEM('o017272, 16'o010605);
`MEM('o017274, 16'o012767);
`MEM('o017276, 16'o021660);
`MEM('o017300, 16'o004664);
`MEM('o017302, 16'o016700);
`MEM('o017304, 16'o004660);
`MEM('o017306, 16'o111000);
`MEM('o017310, 16'o042700);
`MEM('o017312, 16'o177400);
`MEM('o017314, 16'o020027);
`MEM('o017316, 16'o000041);
`MEM('o017320, 16'o001412);
`MEM('o017322, 16'o020027);
`MEM('o017324, 16'o000041);
`MEM('o017326, 16'o003073);
`MEM('o017330, 16'o020027);
`MEM('o017332, 16'o000037);
`MEM('o017334, 16'o001426);
`MEM('o017336, 16'o020027);
`MEM('o017340, 16'o000040);
`MEM('o017342, 16'o001455);
`MEM('o017344, 16'o000464);
`MEM('o017346, 16'o016700);
`MEM('o017350, 16'o004614);
`MEM('o017352, 16'o005200);
`MEM('o017354, 16'o010067);
`MEM('o017356, 16'o004606);
`MEM('o017360, 16'o016700);
`MEM('o017362, 16'o004602);
`MEM('o017364, 16'o111000);
`MEM('o017366, 16'o120027);
`MEM('o017370, 16'o000045);
`MEM('o017372, 16'o001003);
`MEM('o017374, 16'o004767);
`MEM('o017376, 16'o177506);
`MEM('o017400, 16'o000451);
`MEM('o017402, 16'o112767);
`MEM('o017404, 16'o000024);
`MEM('o017406, 16'o001240);
`MEM('o017410, 16'o000445);
`MEM('o017412, 16'o016700);
`MEM('o017414, 16'o004550);
`MEM('o017416, 16'o005200);
`MEM('o017420, 16'o010067);
`MEM('o017422, 16'o004542);
`MEM('o017424, 16'o016700);
`MEM('o017426, 16'o004536);
`MEM('o017430, 16'o111000);
`MEM('o017432, 16'o120027);
`MEM('o017434, 16'o000045);
`MEM('o017436, 16'o001410);
`MEM('o017440, 16'o016700);
`MEM('o017442, 16'o004522);
`MEM('o017444, 16'o062700);
`MEM('o017446, 16'o000003);
`MEM('o017450, 16'o111000);
`MEM('o017452, 16'o120027);
`MEM('o017454, 16'o000045);
`MEM('o017456, 16'o001003);
`MEM('o017460, 16'o004767);
`MEM('o017462, 16'o177074);
`MEM('o017464, 16'o000417);
`MEM('o017466, 16'o112767);
`MEM('o017470, 16'o000024);
`MEM('o017472, 16'o001154);
`MEM('o017474, 16'o000413);
`MEM('o017476, 16'o016700);
`MEM('o017500, 16'o004464);
`MEM('o017502, 16'o005200);
`MEM('o017504, 16'o010067);
`MEM('o017506, 16'o004456);
`MEM('o017510, 16'o004767);
`MEM('o017512, 16'o176726);
`MEM('o017514, 16'o000403);
`MEM('o017516, 16'o004767);
`MEM('o017520, 16'o174164);
`MEM('o017522, 16'o000240);
`MEM('o017524, 16'o000240);
`MEM('o017526, 16'o012605);
`MEM('o017530, 16'o000207);
`MEM('o017532, 16'o010546);
`MEM('o017534, 16'o010605);
`MEM('o017536, 16'o116700);
`MEM('o017540, 16'o001106);
`MEM('o017542, 16'o105700);
`MEM('o017544, 16'o001503);
`MEM('o017546, 16'o016700);
`MEM('o017550, 16'o004414);
`MEM('o017552, 16'o020027);
`MEM('o017554, 16'o022164);
`MEM('o017556, 16'o103460);
`MEM('o017560, 16'o016701);
`MEM('o017562, 16'o004402);
`MEM('o017564, 16'o012700);
`MEM('o017566, 16'o024164);
`MEM('o017570, 16'o020100);
`MEM('o017572, 16'o103052);
`MEM('o017574, 16'o016700);
`MEM('o017576, 16'o004364);
`MEM('o017600, 16'o111000);
`MEM('o017602, 16'o105700);
`MEM('o017604, 16'o001445);
`MEM('o017606, 16'o004767);
`MEM('o017610, 16'o161326);
`MEM('o017612, 16'o012746);
`MEM('o017614, 16'o024452);
`MEM('o017616, 16'o004767);
`MEM('o017620, 16'o161742);
`MEM('o017622, 16'o062706);
`MEM('o017624, 16'o000002);
`MEM('o017626, 16'o016700);
`MEM('o017630, 16'o004332);
`MEM('o017632, 16'o010046);
`MEM('o017634, 16'o004767);
`MEM('o017636, 16'o165624);
`MEM('o017640, 16'o062706);
`MEM('o017642, 16'o000002);
`MEM('o017644, 16'o005046);
`MEM('o017646, 16'o010046);
`MEM('o017650, 16'o004767);
`MEM('o017652, 16'o162360);
`MEM('o017654, 16'o062706);
`MEM('o017656, 16'o000004);
`MEM('o017660, 16'o012746);
`MEM('o017662, 16'o000040);
`MEM('o017664, 16'o004767);
`MEM('o017666, 16'o161120);
`MEM('o017670, 16'o062706);
`MEM('o017672, 16'o000002);
`MEM('o017674, 16'o016700);
`MEM('o017676, 16'o004264);
`MEM('o017700, 16'o062700);
`MEM('o017702, 16'o000003);
`MEM('o017704, 16'o010046);
`MEM('o017706, 16'o004767);
`MEM('o017710, 16'o166544);
`MEM('o017712, 16'o062706);
`MEM('o017714, 16'o000002);
`MEM('o017716, 16'o000416);
`MEM('o017720, 16'o004767);
`MEM('o017722, 16'o161214);
`MEM('o017724, 16'o012746);
`MEM('o017726, 16'o024460);
`MEM('o017730, 16'o004767);
`MEM('o017732, 16'o161630);
`MEM('o017734, 16'o062706);
`MEM('o017736, 16'o000002);
`MEM('o017740, 16'o012746);
`MEM('o017742, 16'o021540);
`MEM('o017744, 16'o004767);
`MEM('o017746, 16'o161614);
`MEM('o017750, 16'o062706);
`MEM('o017752, 16'o000002);
`MEM('o017754, 16'o004767);
`MEM('o017756, 16'o161160);
`MEM('o017760, 16'o116700);
`MEM('o017762, 16'o000664);
`MEM('o017764, 16'o042700);
`MEM('o017766, 16'o177400);
`MEM('o017770, 16'o006300);
`MEM('o017772, 16'o062700);
`MEM('o017774, 16'o021462);
`MEM('o017776, 16'o011000);
`MEM('o020000, 16'o010046);
`MEM('o020002, 16'o004767);
`MEM('o020004, 16'o161556);
`MEM('o020006, 16'o062706);
`MEM('o020010, 16'o000002);
`MEM('o020012, 16'o004767);
`MEM('o020014, 16'o161122);
`MEM('o020016, 16'o105067);
`MEM('o020020, 16'o000626);
`MEM('o020022, 16'o000240);
`MEM('o020024, 16'o012605);
`MEM('o020026, 16'o000207);
`MEM('o020030, 16'o010546);
`MEM('o020032, 16'o010605);
`MEM('o020034, 16'o062706);
`MEM('o020036, 16'o177776);
`MEM('o020040, 16'o004767);
`MEM('o020042, 16'o177042);
`MEM('o020044, 16'o004767);
`MEM('o020046, 16'o161070);
`MEM('o020050, 16'o012746);
`MEM('o020052, 16'o024473);
`MEM('o020054, 16'o004767);
`MEM('o020056, 16'o161504);
`MEM('o020060, 16'o062706);
`MEM('o020062, 16'o000002);
`MEM('o020064, 16'o004767);
`MEM('o020066, 16'o161050);
`MEM('o020070, 16'o012746);
`MEM('o020072, 16'o024520);
`MEM('o020074, 16'o004767);
`MEM('o020076, 16'o161464);
`MEM('o020100, 16'o062706);
`MEM('o020102, 16'o000002);
`MEM('o020104, 16'o012746);
`MEM('o020106, 16'o024527);
`MEM('o020110, 16'o004767);
`MEM('o020112, 16'o161450);
`MEM('o020114, 16'o062706);
`MEM('o020116, 16'o000002);
`MEM('o020120, 16'o004767);
`MEM('o020122, 16'o161014);
`MEM('o020124, 16'o004767);
`MEM('o020126, 16'o177402);
`MEM('o020130, 16'o012746);
`MEM('o020132, 16'o000076);
`MEM('o020134, 16'o004767);
`MEM('o020136, 16'o160650);
`MEM('o020140, 16'o062706);
`MEM('o020142, 16'o000002);
`MEM('o020144, 16'o004767);
`MEM('o020146, 16'o161474);
`MEM('o020150, 16'o004767);
`MEM('o020152, 16'o163142);
`MEM('o020154, 16'o110065);
`MEM('o020156, 16'o177777);
`MEM('o020160, 16'o116700);
`MEM('o020162, 16'o000464);
`MEM('o020164, 16'o105700);
`MEM('o020166, 16'o001403);
`MEM('o020170, 16'o004767);
`MEM('o020172, 16'o177336);
`MEM('o020174, 16'o000427);
`MEM('o020176, 16'o116700);
`MEM('o020200, 16'o001456);
`MEM('o020202, 16'o120027);
`MEM('o020204, 16'o000042);
`MEM('o020206, 16'o001014);
`MEM('o020210, 16'o116567);
`MEM('o020212, 16'o177777);
`MEM('o020214, 16'o001442);
`MEM('o020216, 16'o004767);
`MEM('o020220, 16'o165434);
`MEM('o020222, 16'o116700);
`MEM('o020224, 16'o000422);
`MEM('o020226, 16'o105700);
`MEM('o020230, 16'o001410);
`MEM('o020232, 16'o004767);
`MEM('o020234, 16'o177274);
`MEM('o020236, 16'o000405);
`MEM('o020240, 16'o004767);
`MEM('o020242, 16'o177024);
`MEM('o020244, 16'o004767);
`MEM('o020246, 16'o177262);
`MEM('o020250, 16'o000727);
`MEM('o020252, 16'o000240);
`MEM('o020254, 16'o000725);
`MEM('o020256, 16'o000000);
`MEM('o020260, 16'o000000);
`MEM('o020262, 16'o000000);
`MEM('o020264, 16'o000000);
`MEM('o020266, 16'o000000);
`MEM('o020270, 16'o000000);
`MEM('o020272, 16'o000000);
`MEM('o020274, 16'o000000);
`MEM('o020276, 16'o000000);
`MEM('o020300, 16'o177560);
`MEM('o020302, 16'o177562);
`MEM('o020304, 16'o177564);
`MEM('o020306, 16'o177566);
`MEM('o020310, 16'o047507);
`MEM('o020312, 16'o047524);
`MEM('o020314, 16'o043400);
`MEM('o020316, 16'o051517);
`MEM('o020320, 16'o041125);
`MEM('o020322, 16'o051000);
`MEM('o020324, 16'o052105);
`MEM('o020326, 16'o051125);
`MEM('o020330, 16'o000116);
`MEM('o020332, 16'o047506);
`MEM('o020334, 16'o000122);
`MEM('o020336, 16'o047524);
`MEM('o020340, 16'o051400);
`MEM('o020342, 16'o042524);
`MEM('o020344, 16'o000120);
`MEM('o020346, 16'o042516);
`MEM('o020350, 16'o052130);
`MEM('o020352, 16'o044400);
`MEM('o020354, 16'o000106);
`MEM('o020356, 16'o042522);
`MEM('o020360, 16'o000115);
`MEM('o020362, 16'o052123);
`MEM('o020364, 16'o050117);
`MEM('o020366, 16'o044400);
`MEM('o020370, 16'o050116);
`MEM('o020372, 16'o052125);
`MEM('o020374, 16'o050000);
`MEM('o020376, 16'o044522);
`MEM('o020400, 16'o052116);
`MEM('o020402, 16'o046000);
`MEM('o020404, 16'o052105);
`MEM('o020406, 16'o026000);
`MEM('o020410, 16'o035400);
`MEM('o020412, 16'o026400);
`MEM('o020414, 16'o025400);
`MEM('o020416, 16'o025000);
`MEM('o020420, 16'o027400);
`MEM('o020422, 16'o024000);
`MEM('o020424, 16'o024400);
`MEM('o020426, 16'o037000);
`MEM('o020430, 16'o000075);
`MEM('o020432, 16'o000043);
`MEM('o020434, 16'o000076);
`MEM('o020436, 16'o000075);
`MEM('o020440, 16'o036474);
`MEM('o020442, 16'o036000);
`MEM('o020444, 16'o040000);
`MEM('o020446, 16'o051000);
`MEM('o020450, 16'o042116);
`MEM('o020452, 16'o040400);
`MEM('o020454, 16'o051502);
`MEM('o020456, 16'o051400);
`MEM('o020460, 16'o055111);
`MEM('o020462, 16'o000105);
`MEM('o020464, 16'o044514);
`MEM('o020466, 16'o052123);
`MEM('o020470, 16'o051000);
`MEM('o020472, 16'o047125);
`MEM('o020474, 16'o047000);
`MEM('o020476, 16'o053505);
`MEM('o020500, 16'o000000);
`MEM('o020502, 16'o020310);
`MEM('o020504, 16'o020315);
`MEM('o020506, 16'o020323);
`MEM('o020510, 16'o020332);
`MEM('o020512, 16'o020336);
`MEM('o020514, 16'o020341);
`MEM('o020516, 16'o020346);
`MEM('o020520, 16'o020353);
`MEM('o020522, 16'o020356);
`MEM('o020524, 16'o020362);
`MEM('o020526, 16'o020367);
`MEM('o020530, 16'o020375);
`MEM('o020532, 16'o020403);
`MEM('o020534, 16'o020407);
`MEM('o020536, 16'o020411);
`MEM('o020540, 16'o020413);
`MEM('o020542, 16'o020415);
`MEM('o020544, 16'o020417);
`MEM('o020546, 16'o020421);
`MEM('o020550, 16'o020423);
`MEM('o020552, 16'o020425);
`MEM('o020554, 16'o020427);
`MEM('o020556, 16'o020432);
`MEM('o020560, 16'o020434);
`MEM('o020562, 16'o020436);
`MEM('o020564, 16'o020440);
`MEM('o020566, 16'o020443);
`MEM('o020570, 16'o020445);
`MEM('o020572, 16'o020447);
`MEM('o020574, 16'o020453);
`MEM('o020576, 16'o020457);
`MEM('o020600, 16'o020464);
`MEM('o020602, 16'o020471);
`MEM('o020604, 16'o020475);
`MEM('o020606, 16'o004402);
`MEM('o020610, 16'o007415);
`MEM('o020612, 16'o010420);
`MEM('o020614, 16'o011422);
`MEM('o020616, 16'o012424);
`MEM('o020620, 16'o013426);
`MEM('o020622, 16'o014430);
`MEM('o020624, 16'o015432);
`MEM('o020626, 16'o016434);
`MEM('o020630, 16'o007436);
`MEM('o020632, 16'o010420);
`MEM('o020634, 16'o011422);
`MEM('o020636, 16'o012424);
`MEM('o020640, 16'o013426);
`MEM('o020642, 16'o014430);
`MEM('o020644, 16'o006432);
`MEM('o020646, 16'o022416);
`MEM('o020650, 16'o047400);
`MEM('o020652, 16'o000113);
`MEM('o020654, 16'o062504);
`MEM('o020656, 16'o064566);
`MEM('o020660, 16'o064563);
`MEM('o020662, 16'o067157);
`MEM('o020664, 16'o061040);
`MEM('o020666, 16'o020171);
`MEM('o020670, 16'o062572);
`MEM('o020672, 16'o067562);
`MEM('o020674, 16'o047400);
`MEM('o020676, 16'o062566);
`MEM('o020700, 16'o063162);
`MEM('o020702, 16'o067554);
`MEM('o020704, 16'o000167);
`MEM('o020706, 16'o072523);
`MEM('o020710, 16'o071542);
`MEM('o020712, 16'o071143);
`MEM('o020714, 16'o070151);
`MEM('o020716, 16'o020164);
`MEM('o020720, 16'o072557);
`MEM('o020722, 16'o020164);
`MEM('o020724, 16'o063157);
`MEM('o020726, 16'o071040);
`MEM('o020730, 16'o067141);
`MEM('o020732, 16'o062547);
`MEM('o020734, 16'o044400);
`MEM('o020736, 16'o067543);
`MEM('o020740, 16'o062544);
`MEM('o020742, 16'o061040);
`MEM('o020744, 16'o063165);
`MEM('o020746, 16'o062546);
`MEM('o020750, 16'o020162);
`MEM('o020752, 16'o072546);
`MEM('o020754, 16'o066154);
`MEM('o020756, 16'o046000);
`MEM('o020760, 16'o071551);
`MEM('o020762, 16'o020164);
`MEM('o020764, 16'o072546);
`MEM('o020766, 16'o066154);
`MEM('o020770, 16'o043400);
`MEM('o020772, 16'o051517);
`MEM('o020774, 16'o041125);
`MEM('o020776, 16'o072040);
`MEM('o021000, 16'o067557);
`MEM('o021002, 16'o066440);
`MEM('o021004, 16'o067141);
`MEM('o021006, 16'o020171);
`MEM('o021010, 16'o062556);
`MEM('o021012, 16'o072163);
`MEM('o021014, 16'o062145);
`MEM('o021016, 16'o051000);
`MEM('o021020, 16'o052105);
`MEM('o021022, 16'o051125);
`MEM('o021024, 16'o020116);
`MEM('o021026, 16'o072163);
`MEM('o021030, 16'o061541);
`MEM('o021032, 16'o020153);
`MEM('o021034, 16'o067165);
`MEM('o021036, 16'o062544);
`MEM('o021040, 16'o063162);
`MEM('o021042, 16'o067554);
`MEM('o021044, 16'o000167);
`MEM('o021046, 16'o047506);
`MEM('o021050, 16'o020122);
`MEM('o021052, 16'o067564);
`MEM('o021054, 16'o020157);
`MEM('o021056, 16'o060555);
`MEM('o021060, 16'o074556);
`MEM('o021062, 16'o067040);
`MEM('o021064, 16'o071545);
`MEM('o021066, 16'o062564);
`MEM('o021070, 16'o000144);
`MEM('o021072, 16'o042516);
`MEM('o021074, 16'o052130);
`MEM('o021076, 16'o073440);
`MEM('o021100, 16'o072151);
`MEM('o021102, 16'o067550);
`MEM('o021104, 16'o072165);
`MEM('o021106, 16'o043040);
`MEM('o021110, 16'o051117);
`MEM('o021112, 16'o047000);
`MEM('o021114, 16'o054105);
`MEM('o021116, 16'o020124);
`MEM('o021120, 16'o064567);
`MEM('o021122, 16'o064164);
`MEM('o021124, 16'o072557);
`MEM('o021126, 16'o020164);
`MEM('o021130, 16'o067543);
`MEM('o021132, 16'o067165);
`MEM('o021134, 16'o062564);
`MEM('o021136, 16'o000162);
`MEM('o021140, 16'o042516);
`MEM('o021142, 16'o052130);
`MEM('o021144, 16'o066440);
`MEM('o021146, 16'o071551);
`MEM('o021150, 16'o060555);
`MEM('o021152, 16'o061564);
`MEM('o021154, 16'o020150);
`MEM('o021156, 16'o047506);
`MEM('o021160, 16'o000122);
`MEM('o021162, 16'o047506);
`MEM('o021164, 16'o020122);
`MEM('o021166, 16'o064567);
`MEM('o021170, 16'o064164);
`MEM('o021172, 16'o072557);
`MEM('o021174, 16'o020164);
`MEM('o021176, 16'o060566);
`MEM('o021200, 16'o064562);
`MEM('o021202, 16'o061141);
`MEM('o021204, 16'o062554);
`MEM('o021206, 16'o043000);
`MEM('o021210, 16'o051117);
`MEM('o021212, 16'o073440);
`MEM('o021214, 16'o072151);
`MEM('o021216, 16'o067550);
`MEM('o021220, 16'o072165);
`MEM('o021222, 16'o052040);
`MEM('o021224, 16'o000117);
`MEM('o021226, 16'o042514);
`MEM('o021230, 16'o020124);
`MEM('o021232, 16'o064567);
`MEM('o021234, 16'o064164);
`MEM('o021236, 16'o072557);
`MEM('o021240, 16'o020164);
`MEM('o021242, 16'o060566);
`MEM('o021244, 16'o064562);
`MEM('o021246, 16'o061141);
`MEM('o021250, 16'o062554);
`MEM('o021252, 16'o044400);
`MEM('o021254, 16'o020106);
`MEM('o021256, 16'o064567);
`MEM('o021260, 16'o064164);
`MEM('o021262, 16'o072557);
`MEM('o021264, 16'o020164);
`MEM('o021266, 16'o067543);
`MEM('o021270, 16'o062156);
`MEM('o021272, 16'o072151);
`MEM('o021274, 16'o067551);
`MEM('o021276, 16'o000156);
`MEM('o021300, 16'o067125);
`MEM('o021302, 16'o062544);
`MEM('o021304, 16'o064546);
`MEM('o021306, 16'o062556);
`MEM('o021310, 16'o020144);
`MEM('o021312, 16'o064554);
`MEM('o021314, 16'o062556);
`MEM('o021316, 16'o067040);
`MEM('o021320, 16'o066565);
`MEM('o021322, 16'o062542);
`MEM('o021324, 16'o000162);
`MEM('o021326, 16'o024047);
`MEM('o021330, 16'o020047);
`MEM('o021332, 16'o071157);
`MEM('o021334, 16'o023440);
`MEM('o021336, 16'o023451);
`MEM('o021340, 16'o062440);
`MEM('o021342, 16'o070170);
`MEM('o021344, 16'o061545);
`MEM('o021346, 16'o062564);
`MEM('o021350, 16'o000144);
`MEM('o021352, 16'o036447);
`MEM('o021354, 16'o020047);
`MEM('o021356, 16'o074145);
`MEM('o021360, 16'o062560);
`MEM('o021362, 16'o072143);
`MEM('o021364, 16'o062145);
`MEM('o021366, 16'o044400);
`MEM('o021370, 16'o066154);
`MEM('o021372, 16'o063545);
`MEM('o021374, 16'o066141);
`MEM('o021376, 16'o061440);
`MEM('o021400, 16'o066557);
`MEM('o021402, 16'o060555);
`MEM('o021404, 16'o062156);
`MEM('o021406, 16'o051400);
`MEM('o021410, 16'o067171);
`MEM('o021412, 16'o060564);
`MEM('o021414, 16'o020170);
`MEM('o021416, 16'o071145);
`MEM('o021420, 16'o067562);
`MEM('o021422, 16'o000162);
`MEM('o021424, 16'o067111);
`MEM('o021426, 16'o062564);
`MEM('o021430, 16'o067162);
`MEM('o021432, 16'o066141);
`MEM('o021434, 16'o062440);
`MEM('o021436, 16'o071162);
`MEM('o021440, 16'o071157);
`MEM('o021442, 16'o040400);
`MEM('o021444, 16'o067542);
`MEM('o021446, 16'o072162);
`MEM('o021450, 16'o061040);
`MEM('o021452, 16'o020171);
`MEM('o021454, 16'o042533);
`MEM('o021456, 16'o041523);
`MEM('o021460, 16'o000135);
`MEM('o021462, 16'o020651);
`MEM('o021464, 16'o020654);
`MEM('o021466, 16'o020675);
`MEM('o021470, 16'o020706);
`MEM('o021472, 16'o020735);
`MEM('o021474, 16'o020757);
`MEM('o021476, 16'o020771);
`MEM('o021500, 16'o021017);
`MEM('o021502, 16'o021046);
`MEM('o021504, 16'o021072);
`MEM('o021506, 16'o021113);
`MEM('o021510, 16'o021140);
`MEM('o021512, 16'o021162);
`MEM('o021514, 16'o021207);
`MEM('o021516, 16'o021226);
`MEM('o021520, 16'o021253);
`MEM('o021522, 16'o021300);
`MEM('o021524, 16'o021326);
`MEM('o021526, 16'o021352);
`MEM('o021530, 16'o021367);
`MEM('o021532, 16'o021407);
`MEM('o021534, 16'o021424);
`MEM('o021536, 16'o021443);
`MEM('o021540, 16'o000000);
`MEM('o021542, 16'o000000);
`MEM('o021544, 16'o000000);
`MEM('o021546, 16'o000000);
`MEM('o021550, 16'o000000);
`MEM('o021552, 16'o000000);
`MEM('o021554, 16'o000000);
`MEM('o021556, 16'o000000);
`MEM('o021560, 16'o000000);
`MEM('o021562, 16'o000000);
`MEM('o021564, 16'o000000);
`MEM('o021566, 16'o000000);
`MEM('o021570, 16'o000000);
`MEM('o021572, 16'o000000);
`MEM('o021574, 16'o000000);
`MEM('o021576, 16'o000000);
`MEM('o021600, 16'o000000);
`MEM('o021602, 16'o000000);
`MEM('o021604, 16'o000000);
`MEM('o021606, 16'o000000);
`MEM('o021610, 16'o000000);
`MEM('o021612, 16'o000000);
`MEM('o021614, 16'o000000);
`MEM('o021616, 16'o000000);
`MEM('o021620, 16'o000000);
`MEM('o021622, 16'o000000);
`MEM('o021624, 16'o000000);
`MEM('o021626, 16'o000000);
`MEM('o021630, 16'o000000);
`MEM('o021632, 16'o000000);
`MEM('o021634, 16'o000000);
`MEM('o021636, 16'o000000);
`MEM('o021640, 16'o000000);
`MEM('o021642, 16'o000000);
`MEM('o021644, 16'o000000);
`MEM('o021646, 16'o000000);
`MEM('o021650, 16'o000000);
`MEM('o021652, 16'o000000);
`MEM('o021654, 16'o000000);
`MEM('o021656, 16'o000000);
`MEM('o021660, 16'o000000);
`MEM('o021662, 16'o000000);
`MEM('o021664, 16'o000000);
`MEM('o021666, 16'o000000);
`MEM('o021670, 16'o000000);
`MEM('o021672, 16'o000000);
`MEM('o021674, 16'o000000);
`MEM('o021676, 16'o000000);
`MEM('o021700, 16'o000000);
`MEM('o021702, 16'o000000);
`MEM('o021704, 16'o000000);
`MEM('o021706, 16'o000000);
`MEM('o021710, 16'o000000);
`MEM('o021712, 16'o000000);
`MEM('o021714, 16'o000000);
`MEM('o021716, 16'o000000);
`MEM('o021720, 16'o000000);
`MEM('o021722, 16'o000000);
`MEM('o021724, 16'o000000);
`MEM('o021726, 16'o000000);
`MEM('o021730, 16'o000000);
`MEM('o021732, 16'o000000);
`MEM('o021734, 16'o000000);
`MEM('o021736, 16'o000000);
`MEM('o021740, 16'o000000);
`MEM('o021742, 16'o000000);
`MEM('o021744, 16'o000000);
`MEM('o021746, 16'o000000);
`MEM('o021750, 16'o000000);
`MEM('o021752, 16'o000000);
`MEM('o021754, 16'o000000);
`MEM('o021756, 16'o000000);
`MEM('o021760, 16'o000000);
`MEM('o021762, 16'o000000);
`MEM('o021764, 16'o000000);
`MEM('o021766, 16'o000000);
`MEM('o021770, 16'o000000);
`MEM('o021772, 16'o000000);
`MEM('o021774, 16'o000000);
`MEM('o021776, 16'o000000);
`MEM('o022000, 16'o000000);
`MEM('o022002, 16'o000000);
`MEM('o022004, 16'o000000);
`MEM('o022006, 16'o000000);
`MEM('o022010, 16'o000000);
`MEM('o022012, 16'o000000);
`MEM('o022014, 16'o000000);
`MEM('o022016, 16'o000000);
`MEM('o022020, 16'o000000);
`MEM('o022022, 16'o000000);
`MEM('o022024, 16'o000000);
`MEM('o022026, 16'o000000);
`MEM('o022030, 16'o000000);
`MEM('o022032, 16'o000000);
`MEM('o022034, 16'o000000);
`MEM('o022036, 16'o000000);
`MEM('o022040, 16'o000000);
`MEM('o022042, 16'o000000);
`MEM('o022044, 16'o000000);
`MEM('o022046, 16'o000000);
`MEM('o022050, 16'o000000);
`MEM('o022052, 16'o000000);
`MEM('o022054, 16'o000000);
`MEM('o022056, 16'o000000);
`MEM('o022060, 16'o000000);
`MEM('o022062, 16'o000000);
`MEM('o022064, 16'o000000);
`MEM('o022066, 16'o000000);
`MEM('o022070, 16'o000000);
`MEM('o022072, 16'o000000);
`MEM('o022074, 16'o000000);
`MEM('o022076, 16'o000000);
`MEM('o022100, 16'o000000);
`MEM('o022102, 16'o000000);
`MEM('o022104, 16'o000000);
`MEM('o022106, 16'o000000);
`MEM('o022110, 16'o000000);
`MEM('o022112, 16'o000000);
`MEM('o022114, 16'o000000);
`MEM('o022116, 16'o000000);
`MEM('o022120, 16'o000000);
`MEM('o022122, 16'o000000);
`MEM('o022124, 16'o000000);
`MEM('o022126, 16'o000000);
`MEM('o022130, 16'o000000);
`MEM('o022132, 16'o000000);
`MEM('o022134, 16'o000000);
`MEM('o022136, 16'o000000);
`MEM('o022140, 16'o000000);
`MEM('o022142, 16'o000000);
`MEM('o022144, 16'o000000);
`MEM('o022146, 16'o000000);
`MEM('o022150, 16'o000000);
`MEM('o022152, 16'o000000);
`MEM('o022154, 16'o000000);
`MEM('o022156, 16'o000000);
`MEM('o022160, 16'o000000);
`MEM('o022162, 16'o000000);
`MEM('o022164, 16'o000000);
`MEM('o022166, 16'o000000);
`MEM('o022170, 16'o000000);
`MEM('o022172, 16'o000000);
`MEM('o022174, 16'o000000);
`MEM('o022176, 16'o000000);
`MEM('o022200, 16'o000000);
`MEM('o022202, 16'o000000);
`MEM('o022204, 16'o000000);
`MEM('o022206, 16'o000000);
`MEM('o022210, 16'o000000);
`MEM('o022212, 16'o000000);
`MEM('o022214, 16'o000000);
`MEM('o022216, 16'o000000);
`MEM('o022220, 16'o000000);
`MEM('o022222, 16'o000000);
`MEM('o022224, 16'o000000);
`MEM('o022226, 16'o000000);
`MEM('o022230, 16'o000000);
`MEM('o022232, 16'o000000);
`MEM('o022234, 16'o000000);
`MEM('o022236, 16'o000000);
`MEM('o022240, 16'o000000);
`MEM('o022242, 16'o000000);
`MEM('o022244, 16'o000000);
`MEM('o022246, 16'o000000);
`MEM('o022250, 16'o000000);
`MEM('o022252, 16'o000000);
`MEM('o022254, 16'o000000);
`MEM('o022256, 16'o000000);
`MEM('o022260, 16'o000000);
`MEM('o022262, 16'o000000);
`MEM('o022264, 16'o000000);
`MEM('o022266, 16'o000000);
`MEM('o022270, 16'o000000);
`MEM('o022272, 16'o000000);
`MEM('o022274, 16'o000000);
`MEM('o022276, 16'o000000);
`MEM('o022300, 16'o000000);
`MEM('o022302, 16'o000000);
`MEM('o022304, 16'o000000);
`MEM('o022306, 16'o000000);
`MEM('o022310, 16'o000000);
`MEM('o022312, 16'o000000);
`MEM('o022314, 16'o000000);
`MEM('o022316, 16'o000000);
`MEM('o022320, 16'o000000);
`MEM('o022322, 16'o000000);
`MEM('o022324, 16'o000000);
`MEM('o022326, 16'o000000);
`MEM('o022330, 16'o000000);
`MEM('o022332, 16'o000000);
`MEM('o022334, 16'o000000);
`MEM('o022336, 16'o000000);
`MEM('o022340, 16'o000000);
`MEM('o022342, 16'o000000);
`MEM('o022344, 16'o000000);
`MEM('o022346, 16'o000000);
`MEM('o022350, 16'o000000);
`MEM('o022352, 16'o000000);
`MEM('o022354, 16'o000000);
`MEM('o022356, 16'o000000);
`MEM('o022360, 16'o000000);
`MEM('o022362, 16'o000000);
`MEM('o022364, 16'o000000);
`MEM('o022366, 16'o000000);
`MEM('o022370, 16'o000000);
`MEM('o022372, 16'o000000);
`MEM('o022374, 16'o000000);
`MEM('o022376, 16'o000000);
`MEM('o022400, 16'o000000);
`MEM('o022402, 16'o000000);
`MEM('o022404, 16'o000000);
`MEM('o022406, 16'o000000);
`MEM('o022410, 16'o000000);
`MEM('o022412, 16'o000000);
`MEM('o022414, 16'o000000);
`MEM('o022416, 16'o000000);
`MEM('o022420, 16'o000000);
`MEM('o022422, 16'o000000);
`MEM('o022424, 16'o000000);
`MEM('o022426, 16'o000000);
`MEM('o022430, 16'o000000);
`MEM('o022432, 16'o000000);
`MEM('o022434, 16'o000000);
`MEM('o022436, 16'o000000);
`MEM('o022440, 16'o000000);
`MEM('o022442, 16'o000000);
`MEM('o022444, 16'o000000);
`MEM('o022446, 16'o000000);
`MEM('o022450, 16'o000000);
`MEM('o022452, 16'o000000);
`MEM('o022454, 16'o000000);
`MEM('o022456, 16'o000000);
`MEM('o022460, 16'o000000);
`MEM('o022462, 16'o000000);
`MEM('o022464, 16'o000000);
`MEM('o022466, 16'o000000);
`MEM('o022470, 16'o000000);
`MEM('o022472, 16'o000000);
`MEM('o022474, 16'o000000);
`MEM('o022476, 16'o000000);
`MEM('o022500, 16'o000000);
`MEM('o022502, 16'o000000);
`MEM('o022504, 16'o000000);
`MEM('o022506, 16'o000000);
`MEM('o022510, 16'o000000);
`MEM('o022512, 16'o000000);
`MEM('o022514, 16'o000000);
`MEM('o022516, 16'o000000);
`MEM('o022520, 16'o000000);
`MEM('o022522, 16'o000000);
`MEM('o022524, 16'o000000);
`MEM('o022526, 16'o000000);
`MEM('o022530, 16'o000000);
`MEM('o022532, 16'o000000);
`MEM('o022534, 16'o000000);
`MEM('o022536, 16'o000000);
`MEM('o022540, 16'o000000);
`MEM('o022542, 16'o000000);
`MEM('o022544, 16'o000000);
`MEM('o022546, 16'o000000);
`MEM('o022550, 16'o000000);
`MEM('o022552, 16'o000000);
`MEM('o022554, 16'o000000);
`MEM('o022556, 16'o000000);
`MEM('o022560, 16'o000000);
`MEM('o022562, 16'o000000);
`MEM('o022564, 16'o000000);
`MEM('o022566, 16'o000000);
`MEM('o022570, 16'o000000);
`MEM('o022572, 16'o000000);
`MEM('o022574, 16'o000000);
`MEM('o022576, 16'o000000);
`MEM('o022600, 16'o000000);
`MEM('o022602, 16'o000000);
`MEM('o022604, 16'o000000);
`MEM('o022606, 16'o000000);
`MEM('o022610, 16'o000000);
`MEM('o022612, 16'o000000);
`MEM('o022614, 16'o000000);
`MEM('o022616, 16'o000000);
`MEM('o022620, 16'o000000);
`MEM('o022622, 16'o000000);
`MEM('o022624, 16'o000000);
`MEM('o022626, 16'o000000);
`MEM('o022630, 16'o000000);
`MEM('o022632, 16'o000000);
`MEM('o022634, 16'o000000);
`MEM('o022636, 16'o000000);
`MEM('o022640, 16'o000000);
`MEM('o022642, 16'o000000);
`MEM('o022644, 16'o000000);
`MEM('o022646, 16'o000000);
`MEM('o022650, 16'o000000);
`MEM('o022652, 16'o000000);
`MEM('o022654, 16'o000000);
`MEM('o022656, 16'o000000);
`MEM('o022660, 16'o000000);
`MEM('o022662, 16'o000000);
`MEM('o022664, 16'o000000);
`MEM('o022666, 16'o000000);
`MEM('o022670, 16'o000000);
`MEM('o022672, 16'o000000);
`MEM('o022674, 16'o000000);
`MEM('o022676, 16'o000000);
`MEM('o022700, 16'o000000);
`MEM('o022702, 16'o000000);
`MEM('o022704, 16'o000000);
`MEM('o022706, 16'o000000);
`MEM('o022710, 16'o000000);
`MEM('o022712, 16'o000000);
`MEM('o022714, 16'o000000);
`MEM('o022716, 16'o000000);
`MEM('o022720, 16'o000000);
`MEM('o022722, 16'o000000);
`MEM('o022724, 16'o000000);
`MEM('o022726, 16'o000000);
`MEM('o022730, 16'o000000);
`MEM('o022732, 16'o000000);
`MEM('o022734, 16'o000000);
`MEM('o022736, 16'o000000);
`MEM('o022740, 16'o000000);
`MEM('o022742, 16'o000000);
`MEM('o022744, 16'o000000);
`MEM('o022746, 16'o000000);
`MEM('o022750, 16'o000000);
`MEM('o022752, 16'o000000);
`MEM('o022754, 16'o000000);
`MEM('o022756, 16'o000000);
`MEM('o022760, 16'o000000);
`MEM('o022762, 16'o000000);
`MEM('o022764, 16'o000000);
`MEM('o022766, 16'o000000);
`MEM('o022770, 16'o000000);
`MEM('o022772, 16'o000000);
`MEM('o022774, 16'o000000);
`MEM('o022776, 16'o000000);
`MEM('o023000, 16'o000000);
`MEM('o023002, 16'o000000);
`MEM('o023004, 16'o000000);
`MEM('o023006, 16'o000000);
`MEM('o023010, 16'o000000);
`MEM('o023012, 16'o000000);
`MEM('o023014, 16'o000000);
`MEM('o023016, 16'o000000);
`MEM('o023020, 16'o000000);
`MEM('o023022, 16'o000000);
`MEM('o023024, 16'o000000);
`MEM('o023026, 16'o000000);
`MEM('o023030, 16'o000000);
`MEM('o023032, 16'o000000);
`MEM('o023034, 16'o000000);
`MEM('o023036, 16'o000000);
`MEM('o023040, 16'o000000);
`MEM('o023042, 16'o000000);
`MEM('o023044, 16'o000000);
`MEM('o023046, 16'o000000);
`MEM('o023050, 16'o000000);
`MEM('o023052, 16'o000000);
`MEM('o023054, 16'o000000);
`MEM('o023056, 16'o000000);
`MEM('o023060, 16'o000000);
`MEM('o023062, 16'o000000);
`MEM('o023064, 16'o000000);
`MEM('o023066, 16'o000000);
`MEM('o023070, 16'o000000);
`MEM('o023072, 16'o000000);
`MEM('o023074, 16'o000000);
`MEM('o023076, 16'o000000);
`MEM('o023100, 16'o000000);
`MEM('o023102, 16'o000000);
`MEM('o023104, 16'o000000);
`MEM('o023106, 16'o000000);
`MEM('o023110, 16'o000000);
`MEM('o023112, 16'o000000);
`MEM('o023114, 16'o000000);
`MEM('o023116, 16'o000000);
`MEM('o023120, 16'o000000);
`MEM('o023122, 16'o000000);
`MEM('o023124, 16'o000000);
`MEM('o023126, 16'o000000);
`MEM('o023130, 16'o000000);
`MEM('o023132, 16'o000000);
`MEM('o023134, 16'o000000);
`MEM('o023136, 16'o000000);
`MEM('o023140, 16'o000000);
`MEM('o023142, 16'o000000);
`MEM('o023144, 16'o000000);
`MEM('o023146, 16'o000000);
`MEM('o023150, 16'o000000);
`MEM('o023152, 16'o000000);
`MEM('o023154, 16'o000000);
`MEM('o023156, 16'o000000);
`MEM('o023160, 16'o000000);
`MEM('o023162, 16'o000000);
`MEM('o023164, 16'o000000);
`MEM('o023166, 16'o000000);
`MEM('o023170, 16'o000000);
`MEM('o023172, 16'o000000);
`MEM('o023174, 16'o000000);
`MEM('o023176, 16'o000000);
`MEM('o023200, 16'o000000);
`MEM('o023202, 16'o000000);
`MEM('o023204, 16'o000000);
`MEM('o023206, 16'o000000);
`MEM('o023210, 16'o000000);
`MEM('o023212, 16'o000000);
`MEM('o023214, 16'o000000);
`MEM('o023216, 16'o000000);
`MEM('o023220, 16'o000000);
`MEM('o023222, 16'o000000);
`MEM('o023224, 16'o000000);
`MEM('o023226, 16'o000000);
`MEM('o023230, 16'o000000);
`MEM('o023232, 16'o000000);
`MEM('o023234, 16'o000000);
`MEM('o023236, 16'o000000);
`MEM('o023240, 16'o000000);
`MEM('o023242, 16'o000000);
`MEM('o023244, 16'o000000);
`MEM('o023246, 16'o000000);
`MEM('o023250, 16'o000000);
`MEM('o023252, 16'o000000);
`MEM('o023254, 16'o000000);
`MEM('o023256, 16'o000000);
`MEM('o023260, 16'o000000);
`MEM('o023262, 16'o000000);
`MEM('o023264, 16'o000000);
`MEM('o023266, 16'o000000);
`MEM('o023270, 16'o000000);
`MEM('o023272, 16'o000000);
`MEM('o023274, 16'o000000);
`MEM('o023276, 16'o000000);
`MEM('o023300, 16'o000000);
`MEM('o023302, 16'o000000);
`MEM('o023304, 16'o000000);
`MEM('o023306, 16'o000000);
`MEM('o023310, 16'o000000);
`MEM('o023312, 16'o000000);
`MEM('o023314, 16'o000000);
`MEM('o023316, 16'o000000);
`MEM('o023320, 16'o000000);
`MEM('o023322, 16'o000000);
`MEM('o023324, 16'o000000);
`MEM('o023326, 16'o000000);
`MEM('o023330, 16'o000000);
`MEM('o023332, 16'o000000);
`MEM('o023334, 16'o000000);
`MEM('o023336, 16'o000000);
`MEM('o023340, 16'o000000);
`MEM('o023342, 16'o000000);
`MEM('o023344, 16'o000000);
`MEM('o023346, 16'o000000);
`MEM('o023350, 16'o000000);
`MEM('o023352, 16'o000000);
`MEM('o023354, 16'o000000);
`MEM('o023356, 16'o000000);
`MEM('o023360, 16'o000000);
`MEM('o023362, 16'o000000);
`MEM('o023364, 16'o000000);
`MEM('o023366, 16'o000000);
`MEM('o023370, 16'o000000);
`MEM('o023372, 16'o000000);
`MEM('o023374, 16'o000000);
`MEM('o023376, 16'o000000);
`MEM('o023400, 16'o000000);
`MEM('o023402, 16'o000000);
`MEM('o023404, 16'o000000);
`MEM('o023406, 16'o000000);
`MEM('o023410, 16'o000000);
`MEM('o023412, 16'o000000);
`MEM('o023414, 16'o000000);
`MEM('o023416, 16'o000000);
`MEM('o023420, 16'o000000);
`MEM('o023422, 16'o000000);
`MEM('o023424, 16'o000000);
`MEM('o023426, 16'o000000);
`MEM('o023430, 16'o000000);
`MEM('o023432, 16'o000000);
`MEM('o023434, 16'o000000);
`MEM('o023436, 16'o000000);
`MEM('o023440, 16'o000000);
`MEM('o023442, 16'o000000);
`MEM('o023444, 16'o000000);
`MEM('o023446, 16'o000000);
`MEM('o023450, 16'o000000);
`MEM('o023452, 16'o000000);
`MEM('o023454, 16'o000000);
`MEM('o023456, 16'o000000);
`MEM('o023460, 16'o000000);
`MEM('o023462, 16'o000000);
`MEM('o023464, 16'o000000);
`MEM('o023466, 16'o000000);
`MEM('o023470, 16'o000000);
`MEM('o023472, 16'o000000);
`MEM('o023474, 16'o000000);
`MEM('o023476, 16'o000000);
`MEM('o023500, 16'o000000);
`MEM('o023502, 16'o000000);
`MEM('o023504, 16'o000000);
`MEM('o023506, 16'o000000);
`MEM('o023510, 16'o000000);
`MEM('o023512, 16'o000000);
`MEM('o023514, 16'o000000);
`MEM('o023516, 16'o000000);
`MEM('o023520, 16'o000000);
`MEM('o023522, 16'o000000);
`MEM('o023524, 16'o000000);
`MEM('o023526, 16'o000000);
`MEM('o023530, 16'o000000);
`MEM('o023532, 16'o000000);
`MEM('o023534, 16'o000000);
`MEM('o023536, 16'o000000);
`MEM('o023540, 16'o000000);
`MEM('o023542, 16'o000000);
`MEM('o023544, 16'o000000);
`MEM('o023546, 16'o000000);
`MEM('o023550, 16'o000000);
`MEM('o023552, 16'o000000);
`MEM('o023554, 16'o000000);
`MEM('o023556, 16'o000000);
`MEM('o023560, 16'o000000);
`MEM('o023562, 16'o000000);
`MEM('o023564, 16'o000000);
`MEM('o023566, 16'o000000);
`MEM('o023570, 16'o000000);
`MEM('o023572, 16'o000000);
`MEM('o023574, 16'o000000);
`MEM('o023576, 16'o000000);
`MEM('o023600, 16'o000000);
`MEM('o023602, 16'o000000);
`MEM('o023604, 16'o000000);
`MEM('o023606, 16'o000000);
`MEM('o023610, 16'o000000);
`MEM('o023612, 16'o000000);
`MEM('o023614, 16'o000000);
`MEM('o023616, 16'o000000);
`MEM('o023620, 16'o000000);
`MEM('o023622, 16'o000000);
`MEM('o023624, 16'o000000);
`MEM('o023626, 16'o000000);
`MEM('o023630, 16'o000000);
`MEM('o023632, 16'o000000);
`MEM('o023634, 16'o000000);
`MEM('o023636, 16'o000000);
`MEM('o023640, 16'o000000);
`MEM('o023642, 16'o000000);
`MEM('o023644, 16'o000000);
`MEM('o023646, 16'o000000);
`MEM('o023650, 16'o000000);
`MEM('o023652, 16'o000000);
`MEM('o023654, 16'o000000);
`MEM('o023656, 16'o000000);
`MEM('o023660, 16'o000000);
`MEM('o023662, 16'o000000);
`MEM('o023664, 16'o000000);
`MEM('o023666, 16'o000000);
`MEM('o023670, 16'o000000);
`MEM('o023672, 16'o000000);
`MEM('o023674, 16'o000000);
`MEM('o023676, 16'o000000);
`MEM('o023700, 16'o000000);
`MEM('o023702, 16'o000000);
`MEM('o023704, 16'o000000);
`MEM('o023706, 16'o000000);
`MEM('o023710, 16'o000000);
`MEM('o023712, 16'o000000);
`MEM('o023714, 16'o000000);
`MEM('o023716, 16'o000000);
`MEM('o023720, 16'o000000);
`MEM('o023722, 16'o000000);
`MEM('o023724, 16'o000000);
`MEM('o023726, 16'o000000);
`MEM('o023730, 16'o000000);
`MEM('o023732, 16'o000000);
`MEM('o023734, 16'o000000);
`MEM('o023736, 16'o000000);
`MEM('o023740, 16'o000000);
`MEM('o023742, 16'o000000);
`MEM('o023744, 16'o000000);
`MEM('o023746, 16'o000000);
`MEM('o023750, 16'o000000);
`MEM('o023752, 16'o000000);
`MEM('o023754, 16'o000000);
`MEM('o023756, 16'o000000);
`MEM('o023760, 16'o000000);
`MEM('o023762, 16'o000000);
`MEM('o023764, 16'o000000);
`MEM('o023766, 16'o000000);
`MEM('o023770, 16'o000000);
`MEM('o023772, 16'o000000);
`MEM('o023774, 16'o000000);
`MEM('o023776, 16'o000000);
`MEM('o024000, 16'o000000);
`MEM('o024002, 16'o000000);
`MEM('o024004, 16'o000000);
`MEM('o024006, 16'o000000);
`MEM('o024010, 16'o000000);
`MEM('o024012, 16'o000000);
`MEM('o024014, 16'o000000);
`MEM('o024016, 16'o000000);
`MEM('o024020, 16'o000000);
`MEM('o024022, 16'o000000);
`MEM('o024024, 16'o000000);
`MEM('o024026, 16'o000000);
`MEM('o024030, 16'o000000);
`MEM('o024032, 16'o000000);
`MEM('o024034, 16'o000000);
`MEM('o024036, 16'o000000);
`MEM('o024040, 16'o000000);
`MEM('o024042, 16'o000000);
`MEM('o024044, 16'o000000);
`MEM('o024046, 16'o000000);
`MEM('o024050, 16'o000000);
`MEM('o024052, 16'o000000);
`MEM('o024054, 16'o000000);
`MEM('o024056, 16'o000000);
`MEM('o024060, 16'o000000);
`MEM('o024062, 16'o000000);
`MEM('o024064, 16'o000000);
`MEM('o024066, 16'o000000);
`MEM('o024070, 16'o000000);
`MEM('o024072, 16'o000000);
`MEM('o024074, 16'o000000);
`MEM('o024076, 16'o000000);
`MEM('o024100, 16'o000000);
`MEM('o024102, 16'o000000);
`MEM('o024104, 16'o000000);
`MEM('o024106, 16'o000000);
`MEM('o024110, 16'o000000);
`MEM('o024112, 16'o000000);
`MEM('o024114, 16'o000000);
`MEM('o024116, 16'o000000);
`MEM('o024120, 16'o000000);
`MEM('o024122, 16'o000000);
`MEM('o024124, 16'o000000);
`MEM('o024126, 16'o000000);
`MEM('o024130, 16'o000000);
`MEM('o024132, 16'o000000);
`MEM('o024134, 16'o000000);
`MEM('o024136, 16'o000000);
`MEM('o024140, 16'o000000);
`MEM('o024142, 16'o000000);
`MEM('o024144, 16'o000000);
`MEM('o024146, 16'o000000);
`MEM('o024150, 16'o000000);
`MEM('o024152, 16'o000000);
`MEM('o024154, 16'o000000);
`MEM('o024156, 16'o000000);
`MEM('o024160, 16'o000000);
`MEM('o024162, 16'o000000);
`MEM('o024164, 16'o000000);
`MEM('o024166, 16'o000000);
`MEM('o024170, 16'o000000);
`MEM('o024172, 16'o000000);
`MEM('o024174, 16'o000000);
`MEM('o024176, 16'o000000);
`MEM('o024200, 16'o000000);
`MEM('o024202, 16'o000000);
`MEM('o024204, 16'o000000);
`MEM('o024206, 16'o000000);
`MEM('o024210, 16'o000000);
`MEM('o024212, 16'o000000);
`MEM('o024214, 16'o000000);
`MEM('o024216, 16'o000000);
`MEM('o024220, 16'o000000);
`MEM('o024222, 16'o000000);
`MEM('o024224, 16'o000000);
`MEM('o024226, 16'o000000);
`MEM('o024230, 16'o000000);
`MEM('o024232, 16'o000000);
`MEM('o024234, 16'o000000);
`MEM('o024236, 16'o000000);
`MEM('o024240, 16'o000000);
`MEM('o024242, 16'o000000);
`MEM('o024244, 16'o000000);
`MEM('o024246, 16'o010124);
`MEM('o024250, 16'o010076);
`MEM('o024252, 16'o010502);
`MEM('o024254, 16'o010502);
`MEM('o024256, 16'o010226);
`MEM('o024260, 16'o010502);
`MEM('o024262, 16'o010502);
`MEM('o024264, 16'o010502);
`MEM('o024266, 16'o010502);
`MEM('o024270, 16'o010502);
`MEM('o024272, 16'o010502);
`MEM('o024274, 16'o010502);
`MEM('o024276, 16'o010240);
`MEM('o024300, 16'o010502);
`MEM('o024302, 16'o010332);
`MEM('o024304, 16'o010400);
`MEM('o024306, 16'o010502);
`MEM('o024310, 16'o010502);
`MEM('o024312, 16'o010502);
`MEM('o024314, 16'o010002);
`MEM('o024316, 16'o010156);
`MEM('o024320, 16'o011620);
`MEM('o024322, 16'o011336);
`MEM('o024324, 16'o011546);
`MEM('o024326, 16'o011264);
`MEM('o024330, 16'o011474);
`MEM('o024332, 16'o011422);
`MEM('o024334, 16'o024100);
`MEM('o024336, 16'o024400);
`MEM('o024340, 16'o000072);
`MEM('o024342, 16'o014014);
`MEM('o024344, 16'o014154);
`MEM('o024346, 16'o014430);
`MEM('o024350, 16'o014554);
`MEM('o024352, 16'o016332);
`MEM('o024354, 16'o016332);
`MEM('o024356, 16'o015330);
`MEM('o024360, 16'o016016);
`MEM('o024362, 16'o016102);
`MEM('o024364, 16'o016144);
`MEM('o024366, 16'o016264);
`MEM('o024370, 16'o016244);
`MEM('o024372, 16'o016224);
`MEM('o024374, 16'o016332);
`MEM('o024376, 16'o016316);
`MEM('o024400, 16'o016332);
`MEM('o024402, 16'o016332);
`MEM('o024404, 16'o016332);
`MEM('o024406, 16'o016332);
`MEM('o024410, 16'o016332);
`MEM('o024412, 16'o016332);
`MEM('o024414, 16'o016332);
`MEM('o024416, 16'o016332);
`MEM('o024420, 16'o016332);
`MEM('o024422, 16'o016332);
`MEM('o024424, 16'o016332);
`MEM('o024426, 16'o016332);
`MEM('o024430, 16'o016204);
`MEM('o024432, 16'o016332);
`MEM('o024434, 16'o016332);
`MEM('o024436, 16'o016332);
`MEM('o024440, 16'o016304);
`MEM('o024442, 16'o016304);
`MEM('o024444, 16'o016304);
`MEM('o024446, 16'o016332);
`MEM('o024450, 16'o016164);
`MEM('o024452, 16'o044514);
`MEM('o024454, 16'o042516);
`MEM('o024456, 16'o000072);
`MEM('o024460, 16'o047531);
`MEM('o024462, 16'o020125);
`MEM('o024464, 16'o054524);
`MEM('o024466, 16'o042520);
`MEM('o024470, 16'o020072);
`MEM('o024472, 16'o052000);
`MEM('o024474, 16'o054517);
`MEM('o024476, 16'o051517);
`MEM('o024500, 16'o044510);
`MEM('o024502, 16'o044513);
`MEM('o024504, 16'o052040);
`MEM('o024506, 16'o047111);
`MEM('o024510, 16'o020131);
`MEM('o024512, 16'o040502);
`MEM('o024514, 16'o044523);
`MEM('o024516, 16'o000103);
`MEM('o024520, 16'o042120);
`MEM('o024522, 16'o026520);
`MEM('o024524, 16'o030461);
`MEM('o024526, 16'o020000);
`MEM('o024530, 16'o042105);
`MEM('o024532, 16'o052111);
`MEM('o024534, 16'o047511);
`MEM('o024536, 16'o000116);
`MEM('o024540, 16'o000000);
`MEM('o024542, 16'o000000);
`MEM('o024544, 16'o000000);
`MEM('o024546, 16'o000000);
`MEM('o024550, 16'o000000);
`MEM('o024552, 16'o000000);
`MEM('o024554, 16'o000000);
`MEM('o024556, 16'o000000);
`MEM('o024560, 16'o000000);
`MEM('o024562, 16'o000000);
`MEM('o024564, 16'o000000);
`MEM('o024566, 16'o000000);
`MEM('o024570, 16'o000000);
`MEM('o024572, 16'o000000);
`MEM('o024574, 16'o000000);
`MEM('o024576, 16'o000000);
`MEM('o024600, 16'o000000);
`MEM('o024602, 16'o000004);
`MEM('o024604, 16'o000002);
`MEM('o024606, 16'o001000);
`MEM('o024610, 16'o000000);
`MEM('o024612, 16'o000014);
`MEM('o024614, 16'o000042);
`MEM('o024616, 16'o001000);
`MEM('o024620, 16'o000000);
`MEM('o024622, 16'o000022);
`MEM('o024624, 16'o000042);
`MEM('o024626, 16'o020030);
`MEM('o024630, 16'o000000);
`MEM('o024632, 16'o000032);
`MEM('o024634, 16'o000002);
`MEM('o024636, 16'o001010);
`MEM('o024640, 16'o000000);
`MEM('o024642, 16'o000042);
`MEM('o024644, 16'o000043);
`MEM('o024646, 16'o020300);
`MEM('o024650, 16'o000000);
`MEM('o024652, 16'o000054);
`MEM('o024654, 16'o000043);
`MEM('o024656, 16'o020302);
`MEM('o024660, 16'o000000);
`MEM('o024662, 16'o000066);
`MEM('o024664, 16'o000043);
`MEM('o024666, 16'o020304);
`MEM('o024670, 16'o000000);
`MEM('o024672, 16'o000100);
`MEM('o024674, 16'o000043);
`MEM('o024676, 16'o020306);
`MEM('o024700, 16'o000000);
`MEM('o024702, 16'o000112);
`MEM('o024704, 16'o000042);
`MEM('o024706, 16'o001010);
`MEM('o024710, 16'o000000);
`MEM('o024712, 16'o000123);
`MEM('o024714, 16'o000042);
`MEM('o024716, 16'o001050);
`MEM('o024720, 16'o000000);
`MEM('o024722, 16'o000134);
`MEM('o024724, 16'o000042);
`MEM('o024726, 16'o001106);
`MEM('o024730, 16'o000000);
`MEM('o024732, 16'o000145);
`MEM('o024734, 16'o000042);
`MEM('o024736, 16'o001140);
`MEM('o024740, 16'o000000);
`MEM('o024742, 16'o000156);
`MEM('o024744, 16'o000043);
`MEM('o024746, 16'o020502);
`MEM('o024750, 16'o000000);
`MEM('o024752, 16'o000165);
`MEM('o024754, 16'o000043);
`MEM('o024756, 16'o020606);
`MEM('o024760, 16'o000000);
`MEM('o024762, 16'o000174);
`MEM('o024764, 16'o000043);
`MEM('o024766, 16'o020631);
`MEM('o024770, 16'o000000);
`MEM('o024772, 16'o000203);
`MEM('o024774, 16'o000042);
`MEM('o024776, 16'o001202);
`MEM('o025000, 16'o000000);
`MEM('o025002, 16'o000213);
`MEM('o025004, 16'o000043);
`MEM('o025006, 16'o020650);
`MEM('o025010, 16'o000000);
`MEM('o025012, 16'o000220);
`MEM('o025014, 16'o000043);
`MEM('o025016, 16'o021462);
`MEM('o025020, 16'o000000);
`MEM('o025022, 16'o000230);
`MEM('o025024, 16'o000043);
`MEM('o025026, 16'o021540);
`MEM('o025030, 16'o000000);
`MEM('o025032, 16'o000236);
`MEM('o025034, 16'o000043);
`MEM('o025036, 16'o021660);
`MEM('o025040, 16'o000000);
`MEM('o025042, 16'o000244);
`MEM('o025044, 16'o000043);
`MEM('o025046, 16'o022000);
`MEM('o025050, 16'o000000);
`MEM('o025052, 16'o000251);
`MEM('o025054, 16'o000043);
`MEM('o025056, 16'o022064);
`MEM('o025060, 16'o000000);
`MEM('o025062, 16'o000256);
`MEM('o025064, 16'o000043);
`MEM('o025066, 16'o022164);
`MEM('o025070, 16'o000000);
`MEM('o025072, 16'o000267);
`MEM('o025074, 16'o000043);
`MEM('o025076, 16'o024164);
`MEM('o025100, 16'o000000);
`MEM('o025102, 16'o000274);
`MEM('o025104, 16'o000043);
`MEM('o025106, 16'o024166);
`MEM('o025110, 16'o000000);
`MEM('o025112, 16'o000301);
`MEM('o025114, 16'o000043);
`MEM('o025116, 16'o024170);
`MEM('o025120, 16'o000000);
`MEM('o025122, 16'o000307);
`MEM('o025124, 16'o000043);
`MEM('o025126, 16'o024204);
`MEM('o025130, 16'o000000);
`MEM('o025132, 16'o000316);
`MEM('o025134, 16'o000043);
`MEM('o025136, 16'o024206);
`MEM('o025140, 16'o000000);
`MEM('o025142, 16'o000324);
`MEM('o025144, 16'o000043);
`MEM('o025146, 16'o024244);
`MEM('o025150, 16'o000000);
`MEM('o025152, 16'o000333);
`MEM('o025154, 16'o000042);
`MEM('o025156, 16'o001266);
`MEM('o025160, 16'o000000);
`MEM('o025162, 16'o000346);
`MEM('o025164, 16'o000042);
`MEM('o025166, 16'o001334);
`MEM('o025170, 16'o000000);
`MEM('o025172, 16'o000361);
`MEM('o025174, 16'o000042);
`MEM('o025176, 16'o001374);
`MEM('o025200, 16'o000000);
`MEM('o025202, 16'o000374);
`MEM('o025204, 16'o000042);
`MEM('o025206, 16'o001444);
`MEM('o025210, 16'o000000);
`MEM('o025212, 16'o000407);
`MEM('o025214, 16'o000042);
`MEM('o025216, 16'o001504);
`MEM('o025220, 16'o000000);
`MEM('o025222, 16'o000422);
`MEM('o025224, 16'o000042);
`MEM('o025226, 16'o001564);
`MEM('o025230, 16'o000000);
`MEM('o025232, 16'o000432);
`MEM('o025234, 16'o000042);
`MEM('o025236, 16'o001644);
`MEM('o025240, 16'o000000);
`MEM('o025242, 16'o000442);
`MEM('o025244, 16'o000042);
`MEM('o025246, 16'o002234);
`MEM('o025250, 16'o000000);
`MEM('o025252, 16'o000452);
`MEM('o025254, 16'o000042);
`MEM('o025256, 16'o002530);
`MEM('o025260, 16'o000000);
`MEM('o025262, 16'o000462);
`MEM('o025264, 16'o000042);
`MEM('o025266, 16'o003316);
`MEM('o025270, 16'o000000);
`MEM('o025272, 16'o000472);
`MEM('o025274, 16'o000042);
`MEM('o025276, 16'o005400);
`MEM('o025300, 16'o000000);
`MEM('o025302, 16'o000503);
`MEM('o025304, 16'o000042);
`MEM('o025306, 16'o005464);
`MEM('o025310, 16'o000000);
`MEM('o025312, 16'o000516);
`MEM('o025314, 16'o000042);
`MEM('o025316, 16'o005552);
`MEM('o025320, 16'o000000);
`MEM('o025322, 16'o000525);
`MEM('o025324, 16'o000042);
`MEM('o025326, 16'o005656);
`MEM('o025330, 16'o000000);
`MEM('o025332, 16'o000536);
`MEM('o025334, 16'o000042);
`MEM('o025336, 16'o006456);
`MEM('o025340, 16'o000000);
`MEM('o025342, 16'o000547);
`MEM('o025344, 16'o000042);
`MEM('o025346, 16'o007560);
`MEM('o025350, 16'o000000);
`MEM('o025352, 16'o000561);
`MEM('o025354, 16'o000042);
`MEM('o025356, 16'o011162);
`MEM('o025360, 16'o000000);
`MEM('o025362, 16'o000567);
`MEM('o025364, 16'o000042);
`MEM('o025366, 16'o007726);
`MEM('o025370, 16'o000000);
`MEM('o025372, 16'o000577);
`MEM('o025374, 16'o000042);
`MEM('o025376, 16'o010540);
`MEM('o025400, 16'o000000);
`MEM('o025402, 16'o000605);
`MEM('o025404, 16'o000042);
`MEM('o025406, 16'o010774);
`MEM('o025410, 16'o000000);
`MEM('o025412, 16'o000614);
`MEM('o025414, 16'o000042);
`MEM('o025416, 16'o011712);
`MEM('o025420, 16'o000000);
`MEM('o025422, 16'o000624);
`MEM('o025424, 16'o000042);
`MEM('o025426, 16'o012370);
`MEM('o025430, 16'o000000);
`MEM('o025432, 16'o000634);
`MEM('o025434, 16'o000042);
`MEM('o025436, 16'o013250);
`MEM('o025440, 16'o000000);
`MEM('o025442, 16'o000642);
`MEM('o025444, 16'o000042);
`MEM('o025446, 16'o013414);
`MEM('o025450, 16'o000000);
`MEM('o025452, 16'o000652);
`MEM('o025454, 16'o000042);
`MEM('o025456, 16'o013576);
`MEM('o025460, 16'o000000);
`MEM('o025462, 16'o000660);
`MEM('o025464, 16'o000042);
`MEM('o025466, 16'o013706);
`MEM('o025470, 16'o000000);
`MEM('o025472, 16'o000666);
`MEM('o025474, 16'o000042);
`MEM('o025476, 16'o016442);
`MEM('o025500, 16'o000000);
`MEM('o025502, 16'o000674);
`MEM('o025504, 16'o000042);
`MEM('o025506, 16'o016560);
`MEM('o025510, 16'o000000);
`MEM('o025512, 16'o000703);
`MEM('o025514, 16'o000042);
`MEM('o025516, 16'o017106);
`MEM('o025520, 16'o000000);
`MEM('o025522, 16'o000711);
`MEM('o025524, 16'o000042);
`MEM('o025526, 16'o017270);
`MEM('o025530, 16'o000000);
`MEM('o025532, 16'o000717);
`MEM('o025534, 16'o000042);
`MEM('o025536, 16'o017532);
`MEM('o025540, 16'o000000);
`MEM('o025542, 16'o000726);
`MEM('o025544, 16'o072163);
`MEM('o025546, 16'o071141);
`MEM('o025550, 16'o027164);
`MEM('o025552, 16'o000157);
`MEM('o025554, 16'o072163);
`MEM('o025556, 16'o071141);
`MEM('o025560, 16'o000164);
`MEM('o025562, 16'o061537);
`MEM('o025564, 16'o072163);
`MEM('o025566, 16'o071141);
`MEM('o025570, 16'o000164);
`MEM('o025572, 16'o060542);
`MEM('o025574, 16'o064563);
`MEM('o025576, 16'o027143);
`MEM('o025600, 16'o000157);
`MEM('o025602, 16'o051137);
`MEM('o025604, 16'o043505);
`MEM('o025606, 16'o051137);
`MEM('o025610, 16'o051503);
`MEM('o025612, 16'o000122);
`MEM('o025614, 16'o051137);
`MEM('o025616, 16'o043505);
`MEM('o025620, 16'o051137);
`MEM('o025622, 16'o052502);
`MEM('o025624, 16'o000106);
`MEM('o025626, 16'o051137);
`MEM('o025630, 16'o043505);
`MEM('o025632, 16'o054137);
`MEM('o025634, 16'o051503);
`MEM('o025636, 16'o000122);
`MEM('o025640, 16'o051137);
`MEM('o025642, 16'o043505);
`MEM('o025644, 16'o054137);
`MEM('o025646, 16'o052502);
`MEM('o025650, 16'o000106);
`MEM('o025652, 16'o061537);
`MEM('o025654, 16'o070137);
`MEM('o025656, 16'o072165);
`MEM('o025660, 16'o064143);
`MEM('o025662, 16'o057400);
`MEM('o025664, 16'o057543);
`MEM('o025666, 16'o062547);
`MEM('o025670, 16'o061564);
`MEM('o025672, 16'o000150);
`MEM('o025674, 16'o061537);
`MEM('o025676, 16'o065537);
`MEM('o025700, 16'o064142);
`MEM('o025702, 16'o072151);
`MEM('o025704, 16'o057400);
`MEM('o025706, 16'o062556);
`MEM('o025710, 16'o066167);
`MEM('o025712, 16'o067151);
`MEM('o025714, 16'o000145);
`MEM('o025716, 16'o065537);
`MEM('o025720, 16'o072167);
`MEM('o025722, 16'o066142);
`MEM('o025724, 16'o057400);
`MEM('o025726, 16'o057551);
`MEM('o025730, 16'o071556);
`MEM('o025732, 16'o000141);
`MEM('o025734, 16'o064537);
`MEM('o025736, 16'o067137);
`MEM('o025740, 16'o061163);
`MEM('o025742, 16'o057400);
`MEM('o025744, 16'o071563);
`MEM('o025746, 16'o074564);
`MEM('o025750, 16'o062554);
`MEM('o025752, 16'o057400);
`MEM('o025754, 16'o071145);
`MEM('o025756, 16'o000162);
`MEM('o025760, 16'o062537);
`MEM('o025762, 16'o071162);
`MEM('o025764, 16'o071555);
`MEM('o025766, 16'o000147);
`MEM('o025770, 16'o066137);
`MEM('o025772, 16'o072542);
`MEM('o025774, 16'o000146);
`MEM('o025776, 16'o064537);
`MEM('o026000, 16'o072542);
`MEM('o026002, 16'o000146);
`MEM('o026004, 16'o073137);
`MEM('o026006, 16'o071141);
`MEM('o026010, 16'o057400);
`MEM('o026012, 16'o071141);
`MEM('o026014, 16'o000162);
`MEM('o026016, 16'o066137);
`MEM('o026020, 16'o071551);
`MEM('o026022, 16'o061164);
`MEM('o026024, 16'o063165);
`MEM('o026026, 16'o057400);
`MEM('o026030, 16'o066143);
`MEM('o026032, 16'o000160);
`MEM('o026034, 16'o061537);
`MEM('o026036, 16'o070151);
`MEM('o026040, 16'o057400);
`MEM('o026042, 16'o071547);
`MEM('o026044, 16'o065564);
`MEM('o026046, 16'o057400);
`MEM('o026050, 16'o071547);
`MEM('o026052, 16'o065564);
`MEM('o026054, 16'o000151);
`MEM('o026056, 16'o066137);
`MEM('o026060, 16'o072163);
`MEM('o026062, 16'o000153);
`MEM('o026064, 16'o066137);
`MEM('o026066, 16'o072163);
`MEM('o026070, 16'o064553);
`MEM('o026072, 16'o057400);
`MEM('o026074, 16'o057543);
`MEM('o026076, 16'o067564);
`MEM('o026100, 16'o070165);
`MEM('o026102, 16'o062560);
`MEM('o026104, 16'o000162);
`MEM('o026106, 16'o061537);
`MEM('o026110, 16'o064537);
`MEM('o026112, 16'o070163);
`MEM('o026114, 16'o064562);
`MEM('o026116, 16'o072156);
`MEM('o026120, 16'o057400);
`MEM('o026122, 16'o057543);
`MEM('o026124, 16'o071551);
`MEM('o026126, 16'o070163);
`MEM('o026130, 16'o061541);
`MEM('o026132, 16'o000145);
`MEM('o026134, 16'o061537);
`MEM('o026136, 16'o064537);
`MEM('o026140, 16'o062163);
`MEM('o026142, 16'o063551);
`MEM('o026144, 16'o072151);
`MEM('o026146, 16'o057400);
`MEM('o026150, 16'o057543);
`MEM('o026152, 16'o071551);
`MEM('o026154, 16'o066141);
`MEM('o026156, 16'o064160);
`MEM('o026160, 16'o000141);
`MEM('o026162, 16'o061537);
`MEM('o026164, 16'o070137);
`MEM('o026166, 16'o072165);
`MEM('o026170, 16'o000163);
`MEM('o026172, 16'o061537);
`MEM('o026174, 16'o063537);
`MEM('o026176, 16'o072145);
`MEM('o026200, 16'o000163);
`MEM('o026202, 16'o070137);
`MEM('o026204, 16'o072165);
`MEM('o026206, 16'o072556);
`MEM('o026210, 16'o000155);
`MEM('o026212, 16'o063537);
`MEM('o026214, 16'o072145);
`MEM('o026216, 16'o072556);
`MEM('o026220, 16'o000155);
`MEM('o026222, 16'o072137);
`MEM('o026224, 16'o065557);
`MEM('o026226, 16'o067564);
`MEM('o026230, 16'o000151);
`MEM('o026232, 16'o063537);
`MEM('o026234, 16'o072145);
`MEM('o026236, 16'o064563);
`MEM('o026240, 16'o062572);
`MEM('o026242, 16'o057400);
`MEM('o026244, 16'o062547);
`MEM('o026246, 16'o066164);
`MEM('o026250, 16'o067151);
`MEM('o026252, 16'o067145);
`MEM('o026254, 16'o000157);
`MEM('o026256, 16'o063537);
`MEM('o026260, 16'o072145);
`MEM('o026262, 16'o070154);
`MEM('o026264, 16'o057400);
`MEM('o026266, 16'o067151);
`MEM('o026270, 16'o066163);
`MEM('o026272, 16'o071551);
`MEM('o026274, 16'o000164);
`MEM('o026276, 16'o070137);
`MEM('o026300, 16'o072165);
`MEM('o026302, 16'o064554);
`MEM('o026304, 16'o072163);
`MEM('o026306, 16'o057400);
`MEM('o026310, 16'o062547);
`MEM('o026312, 16'o070164);
`MEM('o026314, 16'o071141);
`MEM('o026316, 16'o066541);
`MEM('o026320, 16'o057400);
`MEM('o026322, 16'o062551);
`MEM('o026324, 16'o070170);
`MEM('o026326, 16'o057400);
`MEM('o026330, 16'o073151);
`MEM('o026332, 16'o066141);
`MEM('o026334, 16'o062565);
`MEM('o026336, 16'o057400);
`MEM('o026340, 16'o066551);
`MEM('o026342, 16'o066165);
`MEM('o026344, 16'o057400);
`MEM('o026346, 16'o070151);
`MEM('o026350, 16'o072554);
`MEM('o026352, 16'o000163);
`MEM('o026354, 16'o064537);
`MEM('o026356, 16'o071160);
`MEM('o026360, 16'o067151);
`MEM('o026362, 16'o000164);
`MEM('o026364, 16'o064537);
`MEM('o026366, 16'o067151);
`MEM('o026370, 16'o072560);
`MEM('o026372, 16'o000164);
`MEM('o026374, 16'o064537);
`MEM('o026376, 16'o060566);
`MEM('o026400, 16'o000162);
`MEM('o026402, 16'o064537);
`MEM('o026404, 16'o071141);
`MEM('o026406, 16'o060562);
`MEM('o026410, 16'o000171);
`MEM('o026412, 16'o064537);
`MEM('o026414, 16'o062554);
`MEM('o026416, 16'o000164);
`MEM('o026420, 16'o064537);
`MEM('o026422, 16'o074145);
`MEM('o026424, 16'o000145);
`MEM('o026426, 16'o064537);
`MEM('o026430, 16'o072562);
`MEM('o026432, 16'o000156);
`MEM('o026434, 16'o064537);
`MEM('o026436, 16'o064554);
`MEM('o026440, 16'o072163);
`MEM('o026442, 16'o057400);
`MEM('o026444, 16'o067151);
`MEM('o026446, 16'o073545);
`MEM('o026450, 16'o057400);
`MEM('o026452, 16'o061551);
`MEM('o026454, 16'o066557);
`MEM('o026456, 16'o057400);
`MEM('o026460, 16'o071145);
`MEM('o026462, 16'o067562);
`MEM('o026464, 16'o000162);
`MEM('o026466, 16'o000000);
end
