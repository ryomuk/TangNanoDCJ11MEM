// rom.v
// to be included from the top module at the comple

`define MEM(x, y) {mem_hi[(x)>>1], mem_lo[(x)>>1]}=y

initial
begin
`MEM('o001000, 16'o012706);
`MEM('o001002, 16'o001000);
`MEM('o001004, 16'o004767);
`MEM('o001006, 16'o000120);
`MEM('o001010, 16'o010546);
`MEM('o001012, 16'o010605);
`MEM('o001014, 16'o000240);
`MEM('o001016, 16'o016700);
`MEM('o001020, 16'o000556);
`MEM('o001022, 16'o011000);
`MEM('o001024, 16'o042700);
`MEM('o001026, 16'o177577);
`MEM('o001030, 16'o005700);
`MEM('o001032, 16'o001771);
`MEM('o001034, 16'o016700);
`MEM('o001036, 16'o000542);
`MEM('o001040, 16'o016510);
`MEM('o001042, 16'o000004);
`MEM('o001044, 16'o000240);
`MEM('o001046, 16'o012605);
`MEM('o001050, 16'o000207);
`MEM('o001052, 16'o010546);
`MEM('o001054, 16'o010605);
`MEM('o001056, 16'o000415);
`MEM('o001060, 16'o016500);
`MEM('o001062, 16'o000004);
`MEM('o001064, 16'o010001);
`MEM('o001066, 16'o005201);
`MEM('o001070, 16'o010165);
`MEM('o001072, 16'o000004);
`MEM('o001074, 16'o111000);
`MEM('o001076, 16'o110000);
`MEM('o001100, 16'o010046);
`MEM('o001102, 16'o004767);
`MEM('o001104, 16'o177702);
`MEM('o001106, 16'o062706);
`MEM('o001110, 16'o000002);
`MEM('o001112, 16'o117500);
`MEM('o001114, 16'o000004);
`MEM('o001116, 16'o105700);
`MEM('o001120, 16'o001357);
`MEM('o001122, 16'o005000);
`MEM('o001124, 16'o012605);
`MEM('o001126, 16'o000207);
`MEM('o001130, 16'o010546);
`MEM('o001132, 16'o174046);
`MEM('o001134, 16'o174146);
`MEM('o001136, 16'o010605);
`MEM('o001140, 16'o062706);
`MEM('o001142, 16'o177722);
`MEM('o001144, 16'o012746);
`MEM('o001146, 16'o001604);
`MEM('o001150, 16'o004767);
`MEM('o001152, 16'o177676);
`MEM('o001154, 16'o062706);
`MEM('o001156, 16'o000002);
`MEM('o001160, 16'o012765);
`MEM('o001162, 16'o177764);
`MEM('o001164, 16'o177772);
`MEM('o001166, 16'o000167);
`MEM('o001170, 16'o000346);
`MEM('o001172, 16'o012765);
`MEM('o001174, 16'o177731);
`MEM('o001176, 16'o177774);
`MEM('o001200, 16'o000543);
`MEM('o001202, 16'o177165);
`MEM('o001204, 16'o177774);
`MEM('o001206, 16'o172467);
`MEM('o001210, 16'o000376);
`MEM('o001212, 16'o171001);
`MEM('o001214, 16'o174065);
`MEM('o001216, 16'o177742);
`MEM('o001220, 16'o177165);
`MEM('o001222, 16'o177772);
`MEM('o001224, 16'o172467);
`MEM('o001226, 16'o000370);
`MEM('o001230, 16'o171001);
`MEM('o001232, 16'o174065);
`MEM('o001234, 16'o177732);
`MEM('o001236, 16'o172465);
`MEM('o001240, 16'o177742);
`MEM('o001242, 16'o174065);
`MEM('o001244, 16'o177762);
`MEM('o001246, 16'o172565);
`MEM('o001250, 16'o177732);
`MEM('o001252, 16'o174165);
`MEM('o001254, 16'o177752);
`MEM('o001256, 16'o005065);
`MEM('o001260, 16'o177776);
`MEM('o001262, 16'o000504);
`MEM('o001264, 16'o172465);
`MEM('o001266, 16'o177762);
`MEM('o001270, 16'o171000);
`MEM('o001272, 16'o172565);
`MEM('o001274, 16'o177752);
`MEM('o001276, 16'o171101);
`MEM('o001300, 16'o173001);
`MEM('o001302, 16'o172565);
`MEM('o001304, 16'o177742);
`MEM('o001306, 16'o172001);
`MEM('o001310, 16'o174065);
`MEM('o001312, 16'o177722);
`MEM('o001314, 16'o172465);
`MEM('o001316, 16'o177762);
`MEM('o001320, 16'o172000);
`MEM('o001322, 16'o171065);
`MEM('o001324, 16'o177752);
`MEM('o001326, 16'o172565);
`MEM('o001330, 16'o177732);
`MEM('o001332, 16'o172001);
`MEM('o001334, 16'o174065);
`MEM('o001336, 16'o177752);
`MEM('o001340, 16'o172465);
`MEM('o001342, 16'o177722);
`MEM('o001344, 16'o174065);
`MEM('o001346, 16'o177762);
`MEM('o001350, 16'o172465);
`MEM('o001352, 16'o177762);
`MEM('o001354, 16'o174001);
`MEM('o001356, 16'o171100);
`MEM('o001360, 16'o172465);
`MEM('o001362, 16'o177752);
`MEM('o001364, 16'o171000);
`MEM('o001366, 16'o172001);
`MEM('o001370, 16'o172527);
`MEM('o001372, 16'o040600);
`MEM('o001374, 16'o173500);
`MEM('o001376, 16'o170000);
`MEM('o001400, 16'o003421);
`MEM('o001402, 16'o026527);
`MEM('o001404, 16'o177776);
`MEM('o001406, 16'o000011);
`MEM('o001410, 16'o003403);
`MEM('o001412, 16'o062765);
`MEM('o001414, 16'o000007);
`MEM('o001416, 16'o177776);
`MEM('o001420, 16'o016500);
`MEM('o001422, 16'o177776);
`MEM('o001424, 16'o062700);
`MEM('o001426, 16'o000060);
`MEM('o001430, 16'o010046);
`MEM('o001432, 16'o004767);
`MEM('o001434, 16'o177352);
`MEM('o001436, 16'o062706);
`MEM('o001440, 16'o000002);
`MEM('o001442, 16'o000420);
`MEM('o001444, 16'o026527);
`MEM('o001446, 16'o177776);
`MEM('o001450, 16'o000017);
`MEM('o001452, 16'o001006);
`MEM('o001454, 16'o012746);
`MEM('o001456, 16'o000040);
`MEM('o001460, 16'o004767);
`MEM('o001462, 16'o177324);
`MEM('o001464, 16'o062706);
`MEM('o001466, 16'o000002);
`MEM('o001470, 16'o005265);
`MEM('o001472, 16'o177776);
`MEM('o001474, 16'o026527);
`MEM('o001476, 16'o177776);
`MEM('o001500, 16'o000017);
`MEM('o001502, 16'o003670);
`MEM('o001504, 16'o005265);
`MEM('o001506, 16'o177774);
`MEM('o001510, 16'o026527);
`MEM('o001512, 16'o177774);
`MEM('o001514, 16'o000047);
`MEM('o001516, 16'o003631);
`MEM('o001520, 16'o012746);
`MEM('o001522, 16'o001604);
`MEM('o001524, 16'o004767);
`MEM('o001526, 16'o177322);
`MEM('o001530, 16'o062706);
`MEM('o001532, 16'o000002);
`MEM('o001534, 16'o005265);
`MEM('o001536, 16'o177772);
`MEM('o001540, 16'o026527);
`MEM('o001542, 16'o177772);
`MEM('o001544, 16'o000014);
`MEM('o001546, 16'o003611);
`MEM('o001550, 16'o000777);
`MEM('o001552, 16'o000000);
`MEM('o001554, 16'o000000);
`MEM('o001556, 16'o000000);
`MEM('o001560, 16'o000000);
`MEM('o001562, 16'o000000);
`MEM('o001564, 16'o000000);
`MEM('o001566, 16'o000000);
`MEM('o001570, 16'o000000);
`MEM('o001572, 16'o000000);
`MEM('o001574, 16'o000000);
`MEM('o001576, 16'o000000);
`MEM('o001600, 16'o177564);
`MEM('o001602, 16'o177566);
`MEM('o001604, 16'o005015);
`MEM('o001606, 16'o000000);
`MEM('o001610, 16'o037073);
`MEM('o001612, 16'o114307);
`MEM('o001614, 16'o161202);
`MEM('o001616, 16'o040270);
`MEM('o001620, 16'o037252);
`MEM('o001622, 16'o124353);
`MEM('o001624, 16'o043064);
`MEM('o001626, 16'o113667);
`MEM('o001630, 16'o000000);
`MEM('o001632, 16'o000000);
`MEM('o001634, 16'o000000);
`MEM('o001636, 16'o000000);
`MEM('o001640, 16'o000000);
`MEM('o001642, 16'o000000);
`MEM('o001644, 16'o000000);
`MEM('o001646, 16'o000000);
`MEM('o001650, 16'o000000);
`MEM('o001652, 16'o000000);
`MEM('o001654, 16'o000000);
`MEM('o001656, 16'o000000);
`MEM('o001660, 16'o000000);
`MEM('o001662, 16'o000000);
`MEM('o001664, 16'o000000);
`MEM('o001666, 16'o000000);
`MEM('o001670, 16'o000000);
`MEM('o001672, 16'o000000);
`MEM('o001674, 16'o000000);
`MEM('o001676, 16'o000000);
`MEM('o001700, 16'o000000);
`MEM('o001702, 16'o000004);
`MEM('o001704, 16'o000002);
`MEM('o001706, 16'o001000);
`MEM('o001710, 16'o000000);
`MEM('o001712, 16'o000014);
`MEM('o001714, 16'o000042);
`MEM('o001716, 16'o001000);
`MEM('o001720, 16'o000000);
`MEM('o001722, 16'o000022);
`MEM('o001724, 16'o000042);
`MEM('o001726, 16'o001130);
`MEM('o001730, 16'o000000);
`MEM('o001732, 16'o000032);
`MEM('o001734, 16'o000002);
`MEM('o001736, 16'o001010);
`MEM('o001740, 16'o000000);
`MEM('o001742, 16'o000045);
`MEM('o001744, 16'o000003);
`MEM('o001746, 16'o001600);
`MEM('o001750, 16'o000000);
`MEM('o001752, 16'o000057);
`MEM('o001754, 16'o000003);
`MEM('o001756, 16'o001602);
`MEM('o001760, 16'o000000);
`MEM('o001762, 16'o000071);
`MEM('o001764, 16'o000042);
`MEM('o001766, 16'o001010);
`MEM('o001770, 16'o000000);
`MEM('o001772, 16'o000102);
`MEM('o001774, 16'o000042);
`MEM('o001776, 16'o001052);
`MEM('o002000, 16'o000000);
`MEM('o002002, 16'o000110);
`MEM('o002004, 16'o072163);
`MEM('o002006, 16'o071141);
`MEM('o002010, 16'o027164);
`MEM('o002012, 16'o000157);
`MEM('o002014, 16'o072163);
`MEM('o002016, 16'o071141);
`MEM('o002020, 16'o000164);
`MEM('o002022, 16'o061537);
`MEM('o002024, 16'o072163);
`MEM('o002026, 16'o071141);
`MEM('o002030, 16'o000164);
`MEM('o002032, 16'o071541);
`MEM('o002034, 16'o064543);
`MEM('o002036, 16'o060551);
`MEM('o002040, 16'o072162);
`MEM('o002042, 16'o067456);
`MEM('o002044, 16'o057400);
`MEM('o002046, 16'o041530);
`MEM('o002050, 16'o051123);
`MEM('o002052, 16'o051137);
`MEM('o002054, 16'o043505);
`MEM('o002056, 16'o057400);
`MEM('o002060, 16'o041130);
`MEM('o002062, 16'o043125);
`MEM('o002064, 16'o051137);
`MEM('o002066, 16'o043505);
`MEM('o002070, 16'o057400);
`MEM('o002072, 16'o072560);
`MEM('o002074, 16'o061564);
`MEM('o002076, 16'o060550);
`MEM('o002100, 16'o000162);
`MEM('o002102, 16'o070137);
`MEM('o002104, 16'o072165);
`MEM('o002106, 16'o000163);
`MEM('o002110, 16'o000000);
end
