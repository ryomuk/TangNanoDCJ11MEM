`define MODULE_NAME Integer_Division_Top
`define SIGNED
`define HAS_REMAINDER
