// rom.v
// to be included from the top module at the comple

`define MEM(x, y) {mem_hi[(x)/2], mem_lo[(x)/2]}=y

initial
begin
`MEM('o000000, 16'o000167);
`MEM('o000002, 16'o003040);
`MEM('o000004, 16'o016146);
`MEM('o000006, 16'o000000);
`MEM('o000010, 16'o000012);
`MEM('o000012, 16'o000000);
`MEM('o000014, 16'o000016);
`MEM('o000016, 16'o000000);
`MEM('o000020, 16'o000022);
`MEM('o000022, 16'o000000);
`MEM('o000024, 16'o000026);
`MEM('o000026, 16'o000000);
`MEM('o000030, 16'o000032);
`MEM('o000032, 16'o000000);
`MEM('o000034, 16'o000100);
`MEM('o000036, 16'o000000);
`MEM('o000040, 16'o000000);
`MEM('o000042, 16'o040407);
`MEM('o000044, 16'o000000);
`MEM('o000046, 16'o000000);
`MEM('o000050, 16'o000056);
`MEM('o000052, 16'o000137);
`MEM('o000054, 16'o000056);
`MEM('o000056, 16'o104465);
`MEM('o000060, 16'o001136);
`MEM('o000062, 16'o000000);
`MEM('o000064, 16'o000066);
`MEM('o000066, 16'o000000);
`MEM('o000070, 16'o000072);
`MEM('o000072, 16'o000000);
`MEM('o000074, 16'o000076);
`MEM('o000076, 16'o000000);
`MEM('o000100, 16'o011666);
`MEM('o000102, 16'o000002);
`MEM('o000104, 16'o162716);
`MEM('o000106, 16'o000002);
`MEM('o000110, 16'o013646);
`MEM('o000112, 16'o006216);
`MEM('o000114, 16'o103404);
`MEM('o000116, 16'o006316);
`MEM('o000120, 16'o062716);
`MEM('o000122, 16'o073654);
`MEM('o000124, 16'o013607);
`MEM('o000126, 16'o042716);
`MEM('o000130, 16'o177600);
`MEM('o000132, 16'o012602);
`MEM('o000134, 16'o020227);
`MEM('o000136, 16'o000100);
`MEM('o000140, 16'o003011);
`MEM('o000142, 16'o005067);
`MEM('o000144, 16'o013526);
`MEM('o000146, 16'o012767);
`MEM('o000150, 16'o000001);
`MEM('o000152, 16'o013524);
`MEM('o000154, 16'o016706);
`MEM('o000156, 16'o013532);
`MEM('o000160, 16'o012746);
`MEM('o000162, 16'o004122);
`MEM('o000164, 16'o010146);
`MEM('o000166, 16'o010201);
`MEM('o000170, 16'o012700);
`MEM('o000172, 16'o000233);
`MEM('o000174, 16'o010146);
`MEM('o000176, 16'o104412);
`MEM('o000200, 16'o104402);
`MEM('o000202, 16'o012700);
`MEM('o000204, 16'o000226);
`MEM('o000206, 16'o104466);
`MEM('o000210, 16'o104404);
`MEM('o000212, 16'o104402);
`MEM('o000214, 16'o005726);
`MEM('o000216, 16'o001001);
`MEM('o000220, 16'o104516);
`MEM('o000222, 16'o012601);
`MEM('o000224, 16'o000207);
`MEM('o000226, 16'o051105);
`MEM('o000230, 16'o047522);
`MEM('o000232, 16'o020122);
`MEM('o000234, 16'o020040);
`MEM('o000236, 16'o020040);
`MEM('o000240, 16'o020040);
`MEM('o000242, 16'o052101);
`MEM('o000244, 16'o046040);
`MEM('o000246, 16'o047111);
`MEM('o000250, 16'o020105);
`MEM('o000252, 16'o000000);
`MEM('o000254, 16'o000476);
`MEM('o000256, 16'o000574);
`MEM('o000260, 16'o002312);
`MEM('o000262, 16'o010074);
`MEM('o000264, 16'o011440);
`MEM('o000266, 16'o011506);
`MEM('o000270, 16'o011566);
`MEM('o000272, 16'o011752);
`MEM('o000274, 16'o012216);
`MEM('o000276, 16'o012442);
`MEM('o000300, 16'o012500);
`MEM('o000302, 16'o012550);
`MEM('o000304, 16'o012776);
`MEM('o000306, 16'o013310);
`MEM('o000310, 16'o013324);
`MEM('o000312, 16'o013166);
`MEM('o000314, 16'o013476);
`MEM('o000316, 16'o013470);
`MEM('o000320, 16'o014646);
`MEM('o000322, 16'o014744);
`MEM('o000324, 16'o014666);
`MEM('o000326, 16'o014536);
`MEM('o000330, 16'o013354);
`MEM('o000332, 16'o014662);
`MEM('o000334, 16'o016016);
`MEM('o000336, 16'o011776);
`MEM('o000340, 16'o012036);
`MEM('o000342, 16'o000606);
`MEM('o000344, 16'o000430);
`MEM('o000346, 16'o001224);
`MEM('o000350, 16'o001656);
`MEM('o000352, 16'o001620);
`MEM('o000354, 16'o000644);
`MEM('o000356, 16'o001646);
`MEM('o000360, 16'o002126);
`MEM('o000362, 16'o002010);
`MEM('o000364, 16'o001236);
`MEM('o000366, 16'o001340);
`MEM('o000370, 16'o001436);
`MEM('o000372, 16'o001256);
`MEM('o000374, 16'o001610);
`MEM('o000376, 16'o001536);
`MEM('o000400, 16'o001772);
`MEM('o000402, 16'o001724);
`MEM('o000404, 16'o002346);
`MEM('o000406, 16'o002144);
`MEM('o000410, 16'o002362);
`MEM('o000412, 16'o004574);
`MEM('o000414, 16'o002400);
`MEM('o000416, 16'o002414);
`MEM('o000420, 16'o006010);
`MEM('o000422, 16'o001302);
`MEM('o000424, 16'o001322);
`MEM('o000426, 16'o017012);
`MEM('o000430, 16'o020227);
`MEM('o000432, 16'o000060);
`MEM('o000434, 16'o002415);
`MEM('o000436, 16'o020227);
`MEM('o000440, 16'o000071);
`MEM('o000442, 16'o003002);
`MEM('o000444, 16'o000264);
`MEM('o000446, 16'o000207);
`MEM('o000450, 16'o020227);
`MEM('o000452, 16'o000101);
`MEM('o000454, 16'o002405);
`MEM('o000456, 16'o020227);
`MEM('o000460, 16'o000132);
`MEM('o000462, 16'o003002);
`MEM('o000464, 16'o000257);
`MEM('o000466, 16'o000207);
`MEM('o000470, 16'o000257);
`MEM('o000472, 16'o000262);
`MEM('o000474, 16'o000207);
`MEM('o000476, 16'o010146);
`MEM('o000500, 16'o012701);
`MEM('o000502, 16'o177564);
`MEM('o000504, 16'o005767);
`MEM('o000506, 16'o013166);
`MEM('o000510, 16'o001403);
`MEM('o000512, 16'o016701);
`MEM('o000514, 16'o013170);
`MEM('o000516, 16'o000416);
`MEM('o000520, 16'o005267);
`MEM('o000522, 16'o013146);
`MEM('o000524, 16'o026727);
`MEM('o000526, 16'o013142);
`MEM('o000530, 16'o000110);
`MEM('o000532, 16'o003405);
`MEM('o000534, 16'o010246);
`MEM('o000536, 16'o010046);
`MEM('o000540, 16'o104402);
`MEM('o000542, 16'o012600);
`MEM('o000544, 16'o012602);
`MEM('o000546, 16'o005767);
`MEM('o000550, 16'o013126);
`MEM('o000552, 16'o001406);
`MEM('o000554, 16'o005267);
`MEM('o000556, 16'o013130);
`MEM('o000560, 16'o105711);
`MEM('o000562, 16'o100374);
`MEM('o000564, 16'o110261);
`MEM('o000566, 16'o000002);
`MEM('o000570, 16'o012601);
`MEM('o000572, 16'o000207);
`MEM('o000574, 16'o012767);
`MEM('o000576, 16'o177776);
`MEM('o000600, 16'o013070);
`MEM('o000602, 16'o012700);
`MEM('o000604, 16'o004103);
`MEM('o000606, 16'o112002);
`MEM('o000610, 16'o001770);
`MEM('o000612, 16'o104400);
`MEM('o000614, 16'o000774);
`MEM('o000616, 16'o005767);
`MEM('o000620, 16'o013052);
`MEM('o000622, 16'o001012);
`MEM('o000624, 16'o022703);
`MEM('o000626, 16'o013540);
`MEM('o000630, 16'o103005);
`MEM('o000632, 16'o012702);
`MEM('o000634, 16'o000134);
`MEM('o000636, 16'o104400);
`MEM('o000640, 16'o005303);
`MEM('o000642, 16'o000402);
`MEM('o000644, 16'o012703);
`MEM('o000646, 16'o013540);
`MEM('o000650, 16'o005767);
`MEM('o000652, 16'o013020);
`MEM('o000654, 16'o001437);
`MEM('o000656, 16'o005067);
`MEM('o000660, 16'o013016);
`MEM('o000662, 16'o016702);
`MEM('o000664, 16'o013016);
`MEM('o000666, 16'o020227);
`MEM('o000670, 16'o177560);
`MEM('o000672, 16'o001002);
`MEM('o000674, 16'o005067);
`MEM('o000676, 16'o176660);
`MEM('o000700, 16'o105212);
`MEM('o000702, 16'o005267);
`MEM('o000704, 16'o013002);
`MEM('o000706, 16'o005712);
`MEM('o000710, 16'o100502);
`MEM('o000712, 16'o105712);
`MEM('o000714, 16'o100372);
`MEM('o000716, 16'o016202);
`MEM('o000720, 16'o000002);
`MEM('o000722, 16'o001752);
`MEM('o000724, 16'o042702);
`MEM('o000726, 16'o177600);
`MEM('o000730, 16'o120227);
`MEM('o000732, 16'o000020);
`MEM('o000734, 16'o001457);
`MEM('o000736, 16'o122702);
`MEM('o000740, 16'o000015);
`MEM('o000742, 16'o001011);
`MEM('o000744, 16'o104402);
`MEM('o000746, 16'o012702);
`MEM('o000750, 16'o000012);
`MEM('o000752, 16'o000417);
`MEM('o000754, 16'o005067);
`MEM('o000756, 16'o176600);
`MEM('o000760, 16'o012702);
`MEM('o000762, 16'o177560);
`MEM('o000764, 16'o000746);
`MEM('o000766, 16'o122702);
`MEM('o000770, 16'o000177);
`MEM('o000772, 16'o001711);
`MEM('o000774, 16'o122702);
`MEM('o000776, 16'o000140);
`MEM('o001000, 16'o003445);
`MEM('o001002, 16'o122702);
`MEM('o001004, 16'o000025);
`MEM('o001006, 16'o001422);
`MEM('o001010, 16'o104400);
`MEM('o001012, 16'o110223);
`MEM('o001014, 16'o120227);
`MEM('o001016, 16'o000012);
`MEM('o001020, 16'o001404);
`MEM('o001022, 16'o020327);
`MEM('o001024, 16'o013657);
`MEM('o001026, 16'o103710);
`MEM('o001030, 16'o104431);
`MEM('o001032, 16'o012701);
`MEM('o001034, 16'o013540);
`MEM('o001036, 16'o012767);
`MEM('o001040, 16'o000001);
`MEM('o001042, 16'o012634);
`MEM('o001044, 16'o052767);
`MEM('o001046, 16'o000100);
`MEM('o001050, 16'o176506);
`MEM('o001052, 16'o000207);
`MEM('o001054, 16'o112702);
`MEM('o001056, 16'o000136);
`MEM('o001060, 16'o104400);
`MEM('o001062, 16'o112702);
`MEM('o001064, 16'o000125);
`MEM('o001066, 16'o104400);
`MEM('o001070, 16'o104402);
`MEM('o001072, 16'o000664);
`MEM('o001074, 16'o012767);
`MEM('o001076, 16'o000100);
`MEM('o001100, 16'o176456);
`MEM('o001102, 16'o005046);
`MEM('o001104, 16'o012746);
`MEM('o001106, 16'o003056);
`MEM('o001110, 16'o010246);
`MEM('o001112, 16'o000423);
`MEM('o001114, 16'o104407);
`MEM('o001116, 16'o005067);
`MEM('o001120, 16'o012552);
`MEM('o001122, 16'o012767);
`MEM('o001124, 16'o000001);
`MEM('o001126, 16'o012550);
`MEM('o001130, 16'o005726);
`MEM('o001132, 16'o000167);
`MEM('o001134, 16'o001754);
`MEM('o001136, 16'o010246);
`MEM('o001140, 16'o116702);
`MEM('o001142, 16'o176416);
`MEM('o001144, 16'o042702);
`MEM('o001146, 16'o177600);
`MEM('o001150, 16'o120227);
`MEM('o001152, 16'o000020);
`MEM('o001154, 16'o001402);
`MEM('o001156, 16'o012602);
`MEM('o001160, 16'o000002);
`MEM('o001162, 16'o016746);
`MEM('o001164, 16'o012512);
`MEM('o001166, 16'o012767);
`MEM('o001170, 16'o000001);
`MEM('o001172, 16'o012504);
`MEM('o001174, 16'o012702);
`MEM('o001176, 16'o000136);
`MEM('o001200, 16'o104400);
`MEM('o001202, 16'o012702);
`MEM('o001204, 16'o000120);
`MEM('o001206, 16'o104400);
`MEM('o001210, 16'o012667);
`MEM('o001212, 16'o012464);
`MEM('o001214, 16'o012767);
`MEM('o001216, 16'o000001);
`MEM('o001220, 16'o012460);
`MEM('o001222, 16'o000755);
`MEM('o001224, 16'o112102);
`MEM('o001226, 16'o122702);
`MEM('o001230, 16'o000040);
`MEM('o001232, 16'o001774);
`MEM('o001234, 16'o000207);
`MEM('o001236, 16'o121127);
`MEM('o001240, 16'o000072);
`MEM('o001242, 16'o001404);
`MEM('o001244, 16'o122127);
`MEM('o001246, 16'o000012);
`MEM('o001250, 16'o001372);
`MEM('o001252, 16'o005301);
`MEM('o001254, 16'o000207);
`MEM('o001256, 16'o005067);
`MEM('o001260, 16'o012406);
`MEM('o001262, 16'o005767);
`MEM('o001264, 16'o012400);
`MEM('o001266, 16'o001404);
`MEM('o001270, 16'o016705);
`MEM('o001272, 16'o012372);
`MEM('o001274, 16'o005067);
`MEM('o001276, 16'o012366);
`MEM('o001300, 16'o000207);
`MEM('o001302, 16'o104512);
`MEM('o001304, 16'o005000);
`MEM('o001306, 16'o104512);
`MEM('o001310, 16'o010500);
`MEM('o001312, 16'o104512);
`MEM('o001314, 16'o104512);
`MEM('o001316, 16'o104512);
`MEM('o001320, 16'o000207);
`MEM('o001322, 16'o010200);
`MEM('o001324, 16'o104512);
`MEM('o001326, 16'o010300);
`MEM('o001330, 16'o104512);
`MEM('o001332, 16'o010400);
`MEM('o001334, 16'o104512);
`MEM('o001336, 16'o000207);
`MEM('o001340, 16'o010446);
`MEM('o001342, 16'o010504);
`MEM('o001344, 16'o062704);
`MEM('o001346, 16'o000024);
`MEM('o001350, 16'o020406);
`MEM('o001352, 16'o103014);
`MEM('o001354, 16'o005767);
`MEM('o001356, 16'o012306);
`MEM('o001360, 16'o001006);
`MEM('o001362, 16'o010567);
`MEM('o001364, 16'o012300);
`MEM('o001366, 16'o005205);
`MEM('o001370, 16'o006205);
`MEM('o001372, 16'o000241);
`MEM('o001374, 16'o006305);
`MEM('o001376, 16'o010025);
`MEM('o001400, 16'o012604);
`MEM('o001402, 16'o000207);
`MEM('o001404, 16'o104401);
`MEM('o001406, 16'o011300);
`MEM('o001410, 16'o041600);
`MEM('o001412, 16'o020004);
`MEM('o001414, 16'o001423);
`MEM('o001416, 16'o042700);
`MEM('o001420, 16'o017777);
`MEM('o001422, 16'o022700);
`MEM('o001424, 16'o040000);
`MEM('o001426, 16'o001022);
`MEM('o001430, 16'o062703);
`MEM('o001432, 16'o000020);
`MEM('o001434, 16'o000406);
`MEM('o001436, 16'o005703);
`MEM('o001440, 16'o001414);
`MEM('o001442, 16'o020506);
`MEM('o001444, 16'o103357);
`MEM('o001446, 16'o010146);
`MEM('o001450, 16'o010046);
`MEM('o001452, 16'o020306);
`MEM('o001454, 16'o103353);
`MEM('o001456, 16'o020305);
`MEM('o001460, 16'o103752);
`MEM('o001462, 16'o005003);
`MEM('o001464, 16'o012600);
`MEM('o001466, 16'o012601);
`MEM('o001470, 16'o005703);
`MEM('o001472, 16'o000207);
`MEM('o001474, 16'o003005);
`MEM('o001476, 16'o062703);
`MEM('o001500, 16'o000002);
`MEM('o001502, 16'o062703);
`MEM('o001504, 16'o000004);
`MEM('o001506, 16'o000761);
`MEM('o001510, 16'o005700);
`MEM('o001512, 16'o001402);
`MEM('o001514, 16'o005723);
`MEM('o001516, 16'o000755);
`MEM('o001520, 16'o116300);
`MEM('o001522, 16'o000002);
`MEM('o001524, 16'o116301);
`MEM('o001526, 16'o000003);
`MEM('o001530, 16'o104522);
`MEM('o001532, 16'o060003);
`MEM('o001534, 16'o000762);
`MEM('o001536, 16'o042700);
`MEM('o001540, 16'o177400);
`MEM('o001542, 16'o042701);
`MEM('o001544, 16'o177400);
`MEM('o001546, 16'o005200);
`MEM('o001550, 16'o005201);
`MEM('o001552, 16'o010446);
`MEM('o001554, 16'o010346);
`MEM('o001556, 16'o104416);
`MEM('o001560, 16'o012603);
`MEM('o001562, 16'o012604);
`MEM('o001564, 16'o005701);
`MEM('o001566, 16'o001006);
`MEM('o001570, 16'o020027);
`MEM('o001572, 16'o022000);
`MEM('o001574, 16'o103003);
`MEM('o001576, 16'o104530);
`MEM('o001600, 16'o000257);
`MEM('o001602, 16'o000207);
`MEM('o001604, 16'o000262);
`MEM('o001606, 16'o000207);
`MEM('o001610, 16'o010301);
`MEM('o001612, 16'o010102);
`MEM('o001614, 16'o060401);
`MEM('o001616, 16'o000404);
`MEM('o001620, 16'o104516);
`MEM('o001622, 16'o010103);
`MEM('o001624, 16'o010102);
`MEM('o001626, 16'o104502);
`MEM('o001630, 16'o020105);
`MEM('o001632, 16'o103002);
`MEM('o001634, 16'o112123);
`MEM('o001636, 16'o000774);
`MEM('o001640, 16'o010305);
`MEM('o001642, 16'o010201);
`MEM('o001644, 16'o000207);
`MEM('o001646, 16'o122127);
`MEM('o001650, 16'o000012);
`MEM('o001652, 16'o001375);
`MEM('o001654, 16'o000207);
`MEM('o001656, 16'o016701);
`MEM('o001660, 16'o012000);
`MEM('o001662, 16'o104502);
`MEM('o001664, 16'o020105);
`MEM('o001666, 16'o103013);
`MEM('o001670, 16'o010046);
`MEM('o001672, 16'o010146);
`MEM('o001674, 16'o104410);
`MEM('o001676, 16'o012601);
`MEM('o001700, 16'o010002);
`MEM('o001702, 16'o012600);
`MEM('o001704, 16'o020002);
`MEM('o001706, 16'o001402);
`MEM('o001710, 16'o003364);
`MEM('o001712, 16'o000257);
`MEM('o001714, 16'o000207);
`MEM('o001716, 16'o000257);
`MEM('o001720, 16'o000262);
`MEM('o001722, 16'o000207);
`MEM('o001724, 16'o104472);
`MEM('o001726, 16'o104470);
`MEM('o001730, 16'o001416);
`MEM('o001732, 16'o102415);
`MEM('o001734, 16'o042702);
`MEM('o001736, 16'o177700);
`MEM('o001740, 16'o010204);
`MEM('o001742, 16'o000304);
`MEM('o001744, 16'o006204);
`MEM('o001746, 16'o006204);
`MEM('o001750, 16'o104472);
`MEM('o001752, 16'o104470);
`MEM('o001754, 16'o001002);
`MEM('o001756, 16'o050204);
`MEM('o001760, 16'o104472);
`MEM('o001762, 16'o000257);
`MEM('o001764, 16'o000207);
`MEM('o001766, 16'o000262);
`MEM('o001770, 16'o000207);
`MEM('o001772, 16'o005700);
`MEM('o001774, 16'o002746);
`MEM('o001776, 16'o020027);
`MEM('o002000, 16'o000377);
`MEM('o002002, 16'o003343);
`MEM('o002004, 16'o000264);
`MEM('o002006, 16'o000207);
`MEM('o002010, 16'o104472);
`MEM('o002012, 16'o104470);
`MEM('o002014, 16'o001015);
`MEM('o002016, 16'o005301);
`MEM('o002020, 16'o104410);
`MEM('o002022, 16'o010046);
`MEM('o002024, 16'o104472);
`MEM('o002026, 16'o022702);
`MEM('o002030, 16'o000054);
`MEM('o002032, 16'o001010);
`MEM('o002034, 16'o104410);
`MEM('o002036, 16'o005700);
`MEM('o002040, 16'o001405);
`MEM('o002042, 16'o010004);
`MEM('o002044, 16'o012603);
`MEM('o002046, 16'o000207);
`MEM('o002050, 16'o005046);
`MEM('o002052, 16'o000765);
`MEM('o002054, 16'o005004);
`MEM('o002056, 16'o000772);
`MEM('o002060, 16'o012767);
`MEM('o002062, 16'o000001);
`MEM('o002064, 16'o011610);
`MEM('o002066, 16'o000167);
`MEM('o002070, 16'o000346);
`MEM('o002072, 16'o012767);
`MEM('o002074, 16'o000001);
`MEM('o002076, 16'o011574);
`MEM('o002100, 16'o016705);
`MEM('o002102, 16'o011556);
`MEM('o002104, 16'o005205);
`MEM('o002106, 16'o005067);
`MEM('o002110, 16'o011554);
`MEM('o002112, 16'o005067);
`MEM('o002114, 16'o011564);
`MEM('o002116, 16'o005067);
`MEM('o002120, 16'o011536);
`MEM('o002122, 16'o000167);
`MEM('o002124, 16'o000634);
`MEM('o002126, 16'o010504);
`MEM('o002130, 16'o060004);
`MEM('o002132, 16'o010603);
`MEM('o002134, 16'o162703);
`MEM('o002136, 16'o000070);
`MEM('o002140, 16'o020304);
`MEM('o002142, 16'o000207);
`MEM('o002144, 16'o010346);
`MEM('o002146, 16'o104536);
`MEM('o002150, 16'o102437);
`MEM('o002152, 16'o121127);
`MEM('o002154, 16'o000054);
`MEM('o002156, 16'o001041);
`MEM('o002160, 16'o004767);
`MEM('o002162, 16'o000102);
`MEM('o002164, 16'o104472);
`MEM('o002166, 16'o010046);
`MEM('o002170, 16'o104536);
`MEM('o002172, 16'o102033);
`MEM('o002174, 16'o104440);
`MEM('o002176, 16'o100432);
`MEM('o002200, 16'o012602);
`MEM('o002202, 16'o017604);
`MEM('o002204, 16'o000000);
`MEM('o002206, 16'o042704);
`MEM('o002210, 16'o177400);
`MEM('o002212, 16'o020004);
`MEM('o002214, 16'o003023);
`MEM('o002216, 16'o010146);
`MEM('o002220, 16'o010201);
`MEM('o002222, 16'o010046);
`MEM('o002224, 16'o010400);
`MEM('o002226, 16'o005200);
`MEM('o002230, 16'o104416);
`MEM('o002232, 16'o062600);
`MEM('o002234, 16'o104530);
`MEM('o002236, 16'o012601);
`MEM('o002240, 16'o061600);
`MEM('o002242, 16'o005720);
`MEM('o002244, 16'o012603);
`MEM('o002246, 16'o000207);
`MEM('o002250, 16'o004767);
`MEM('o002252, 16'o000012);
`MEM('o002254, 16'o010002);
`MEM('o002256, 16'o005000);
`MEM('o002260, 16'o000750);
`MEM('o002262, 16'o104413);
`MEM('o002264, 16'o104415);
`MEM('o002266, 16'o104440);
`MEM('o002270, 16'o100775);
`MEM('o002272, 16'o017604);
`MEM('o002274, 16'o000002);
`MEM('o002276, 16'o000304);
`MEM('o002300, 16'o042704);
`MEM('o002302, 16'o177400);
`MEM('o002304, 16'o020004);
`MEM('o002306, 16'o003366);
`MEM('o002310, 16'o000207);
`MEM('o002312, 16'o162706);
`MEM('o002314, 16'o000010);
`MEM('o002316, 16'o010600);
`MEM('o002320, 16'o016701);
`MEM('o002322, 16'o011334);
`MEM('o002324, 16'o104412);
`MEM('o002326, 16'o010600);
`MEM('o002330, 16'o005720);
`MEM('o002332, 16'o105066);
`MEM('o002334, 16'o000007);
`MEM('o002336, 16'o104466);
`MEM('o002340, 16'o062706);
`MEM('o002342, 16'o000010);
`MEM('o002344, 16'o000207);
`MEM('o002346, 16'o000241);
`MEM('o002350, 16'o006300);
`MEM('o002352, 16'o010046);
`MEM('o002354, 16'o006300);
`MEM('o002356, 16'o062600);
`MEM('o002360, 16'o000207);
`MEM('o002362, 16'o016703);
`MEM('o002364, 16'o011300);
`MEM('o002366, 16'o005203);
`MEM('o002370, 16'o006203);
`MEM('o002372, 16'o000241);
`MEM('o002374, 16'o006303);
`MEM('o002376, 16'o000207);
`MEM('o002400, 16'o104472);
`MEM('o002402, 16'o010204);
`MEM('o002404, 16'o000304);
`MEM('o002406, 16'o104472);
`MEM('o002410, 16'o050204);
`MEM('o002412, 16'o000207);
`MEM('o002414, 16'o010346);
`MEM('o002416, 16'o010246);
`MEM('o002420, 16'o016646);
`MEM('o002422, 16'o000004);
`MEM('o002424, 16'o010466);
`MEM('o002426, 16'o000006);
`MEM('o002430, 16'o020506);
`MEM('o002432, 16'o103001);
`MEM('o002434, 16'o000207);
`MEM('o002436, 16'o104401);
`MEM('o002440, 16'o104516);
`MEM('o002442, 16'o104506);
`MEM('o002444, 16'o010300);
`MEM('o002446, 16'o001060);
`MEM('o002450, 16'o016703);
`MEM('o002452, 16'o011206);
`MEM('o002454, 16'o005704);
`MEM('o002456, 16'o001062);
`MEM('o002460, 16'o010504);
`MEM('o002462, 16'o005767);
`MEM('o002464, 16'o011214);
`MEM('o002466, 16'o001076);
`MEM('o002470, 16'o112302);
`MEM('o002472, 16'o120227);
`MEM('o002474, 16'o000140);
`MEM('o002476, 16'o002421);
`MEM('o002500, 16'o162702);
`MEM('o002502, 16'o000140);
`MEM('o002504, 16'o012700);
`MEM('o002506, 16'o003626);
`MEM('o002510, 16'o010201);
`MEM('o002512, 16'o005301);
`MEM('o002514, 16'o002404);
`MEM('o002516, 16'o122027);
`MEM('o002520, 16'o000044);
`MEM('o002522, 16'o001375);
`MEM('o002524, 16'o000772);
`MEM('o002526, 16'o112002);
`MEM('o002530, 16'o120227);
`MEM('o002532, 16'o000044);
`MEM('o002534, 16'o001752);
`MEM('o002536, 16'o104400);
`MEM('o002540, 16'o000772);
`MEM('o002542, 16'o120227);
`MEM('o002544, 16'o000012);
`MEM('o002546, 16'o001402);
`MEM('o002550, 16'o104400);
`MEM('o002552, 16'o000743);
`MEM('o002554, 16'o104402);
`MEM('o002556, 16'o020304);
`MEM('o002560, 16'o103740);
`MEM('o002562, 16'o005767);
`MEM('o002564, 16'o011110);
`MEM('o002566, 16'o001406);
`MEM('o002570, 16'o005002);
`MEM('o002572, 16'o012701);
`MEM('o002574, 16'o000100);
`MEM('o002576, 16'o104400);
`MEM('o002600, 16'o005301);
`MEM('o002602, 16'o001375);
`MEM('o002604, 16'o000167);
`MEM('o002606, 16'o000276);
`MEM('o002610, 16'o010446);
`MEM('o002612, 16'o104474);
`MEM('o002614, 16'o012604);
`MEM('o002616, 16'o020105);
`MEM('o002620, 16'o101313);
`MEM('o002622, 16'o010103);
`MEM('o002624, 16'o020400);
`MEM('o002626, 16'o003407);
`MEM('o002630, 16'o010400);
`MEM('o002632, 16'o010346);
`MEM('o002634, 16'o104474);
`MEM('o002636, 16'o001006);
`MEM('o002640, 16'o012603);
`MEM('o002642, 16'o020105);
`MEM('o002644, 16'o101305);
`MEM('o002646, 16'o104502);
`MEM('o002650, 16'o010104);
`MEM('o002652, 16'o000703);
`MEM('o002654, 16'o012603);
`MEM('o002656, 16'o020105);
`MEM('o002660, 16'o101277);
`MEM('o002662, 16'o000772);
`MEM('o002664, 16'o000167);
`MEM('o002666, 16'o000166);
`MEM('o002670, 16'o104516);
`MEM('o002672, 16'o104506);
`MEM('o002674, 16'o016701);
`MEM('o002676, 16'o010762);
`MEM('o002700, 16'o005704);
`MEM('o002702, 16'o001001);
`MEM('o002704, 16'o010304);
`MEM('o002706, 16'o010446);
`MEM('o002710, 16'o010346);
`MEM('o002712, 16'o104502);
`MEM('o002714, 16'o020105);
`MEM('o002716, 16'o103012);
`MEM('o002720, 16'o010146);
`MEM('o002722, 16'o104410);
`MEM('o002724, 16'o012601);
`MEM('o002726, 16'o020016);
`MEM('o002730, 16'o002770);
`MEM('o002732, 16'o020066);
`MEM('o002734, 16'o000002);
`MEM('o002736, 16'o003002);
`MEM('o002740, 16'o104476);
`MEM('o002742, 16'o000764);
`MEM('o002744, 16'o022626);
`MEM('o002746, 16'o000461);
`MEM('o002750, 16'o104516);
`MEM('o002752, 16'o104474);
`MEM('o002754, 16'o001013);
`MEM('o002756, 16'o104476);
`MEM('o002760, 16'o000411);
`MEM('o002762, 16'o004767);
`MEM('o002764, 16'o176236);
`MEM('o002766, 16'o122702);
`MEM('o002770, 16'o000072);
`MEM('o002772, 16'o001520);
`MEM('o002774, 16'o122702);
`MEM('o002776, 16'o000012);
`MEM('o003000, 16'o001401);
`MEM('o003002, 16'o104407);
`MEM('o003004, 16'o005767);
`MEM('o003006, 16'o010654);
`MEM('o003010, 16'o001445);
`MEM('o003012, 16'o005767);
`MEM('o003014, 16'o010650);
`MEM('o003016, 16'o001403);
`MEM('o003020, 16'o020167);
`MEM('o003022, 16'o010642);
`MEM('o003024, 16'o000401);
`MEM('o003026, 16'o020105);
`MEM('o003030, 16'o103114);
`MEM('o003032, 16'o004767);
`MEM('o003034, 16'o006402);
`MEM('o003036, 16'o010067);
`MEM('o003040, 16'o010616);
`MEM('o003042, 16'o000474);
`MEM('o003044, 16'o016705);
`MEM('o003046, 16'o010612);
`MEM('o003050, 16'o005205);
`MEM('o003052, 16'o005067);
`MEM('o003054, 16'o010610);
`MEM('o003056, 16'o016706);
`MEM('o003060, 16'o010630);
`MEM('o003062, 16'o005067);
`MEM('o003064, 16'o010606);
`MEM('o003066, 16'o005067);
`MEM('o003070, 16'o010610);
`MEM('o003072, 16'o005067);
`MEM('o003074, 16'o010562);
`MEM('o003076, 16'o012767);
`MEM('o003100, 16'o000001);
`MEM('o003102, 16'o010574);
`MEM('o003104, 16'o104402);
`MEM('o003106, 16'o005067);
`MEM('o003110, 16'o010564);
`MEM('o003112, 16'o005067);
`MEM('o003114, 16'o010546);
`MEM('o003116, 16'o012700);
`MEM('o003120, 16'o004076);
`MEM('o003122, 16'o104466);
`MEM('o003124, 16'o005067);
`MEM('o003126, 16'o010552);
`MEM('o003130, 16'o104500);
`MEM('o003132, 16'o104472);
`MEM('o003134, 16'o020227);
`MEM('o003136, 16'o000012);
`MEM('o003140, 16'o001771);
`MEM('o003142, 16'o012701);
`MEM('o003144, 16'o013540);
`MEM('o003146, 16'o104410);
`MEM('o003150, 16'o121127);
`MEM('o003152, 16'o000012);
`MEM('o003154, 16'o001675);
`MEM('o003156, 16'o010103);
`MEM('o003160, 16'o012700);
`MEM('o003162, 16'o003626);
`MEM('o003164, 16'o005002);
`MEM('o003166, 16'o122327);
`MEM('o003170, 16'o000040);
`MEM('o003172, 16'o001775);
`MEM('o003174, 16'o124320);
`MEM('o003176, 16'o001005);
`MEM('o003200, 16'o005203);
`MEM('o003202, 16'o121027);
`MEM('o003204, 16'o000044);
`MEM('o003206, 16'o001430);
`MEM('o003210, 16'o000766);
`MEM('o003212, 16'o122027);
`MEM('o003214, 16'o000044);
`MEM('o003216, 16'o001375);
`MEM('o003220, 16'o121027);
`MEM('o003222, 16'o000044);
`MEM('o003224, 16'o001420);
`MEM('o003226, 16'o010103);
`MEM('o003230, 16'o005202);
`MEM('o003232, 16'o000755);
`MEM('o003234, 16'o005767);
`MEM('o003236, 16'o010442);
`MEM('o003240, 16'o001306);
`MEM('o003242, 16'o004767);
`MEM('o003244, 16'o175756);
`MEM('o003246, 16'o162702);
`MEM('o003250, 16'o000140);
`MEM('o003252, 16'o100405);
`MEM('o003254, 16'o006302);
`MEM('o003256, 16'o000172);
`MEM('o003260, 16'o004020);
`MEM('o003262, 16'o000167);
`MEM('o003264, 16'o000620);
`MEM('o003266, 16'o104403);
`MEM('o003270, 16'o062702);
`MEM('o003272, 16'o000140);
`MEM('o003274, 16'o110221);
`MEM('o003276, 16'o010104);
`MEM('o003300, 16'o111321);
`MEM('o003302, 16'o122327);
`MEM('o003304, 16'o000012);
`MEM('o003306, 16'o001374);
`MEM('o003310, 16'o120227);
`MEM('o003312, 16'o000143);
`MEM('o003314, 16'o001465);
`MEM('o003316, 16'o020227);
`MEM('o003320, 16'o000155);
`MEM('o003322, 16'o001035);
`MEM('o003324, 16'o010401);
`MEM('o003326, 16'o104472);
`MEM('o003330, 16'o120227);
`MEM('o003332, 16'o000124);
`MEM('o003334, 16'o001022);
`MEM('o003336, 16'o104472);
`MEM('o003340, 16'o120227);
`MEM('o003342, 16'o000110);
`MEM('o003344, 16'o001016);
`MEM('o003346, 16'o104472);
`MEM('o003350, 16'o120227);
`MEM('o003352, 16'o000105);
`MEM('o003354, 16'o001012);
`MEM('o003356, 16'o104472);
`MEM('o003360, 16'o120227);
`MEM('o003362, 16'o000116);
`MEM('o003364, 16'o001006);
`MEM('o003366, 16'o104472);
`MEM('o003370, 16'o005301);
`MEM('o003372, 16'o010104);
`MEM('o003374, 16'o104470);
`MEM('o003376, 16'o001407);
`MEM('o003400, 16'o000666);
`MEM('o003402, 16'o120227);
`MEM('o003404, 16'o000012);
`MEM('o003406, 16'o001430);
`MEM('o003410, 16'o120227);
`MEM('o003412, 16'o000072);
`MEM('o003414, 16'o001344);
`MEM('o003416, 16'o010401);
`MEM('o003420, 16'o121127);
`MEM('o003422, 16'o000042);
`MEM('o003424, 16'o001410);
`MEM('o003426, 16'o122127);
`MEM('o003430, 16'o000072);
`MEM('o003432, 16'o001755);
`MEM('o003434, 16'o124127);
`MEM('o003436, 16'o000012);
`MEM('o003440, 16'o001412);
`MEM('o003442, 16'o005201);
`MEM('o003444, 16'o000765);
`MEM('o003446, 16'o005201);
`MEM('o003450, 16'o121127);
`MEM('o003452, 16'o000042);
`MEM('o003454, 16'o001772);
`MEM('o003456, 16'o121127);
`MEM('o003460, 16'o000012);
`MEM('o003462, 16'o001371);
`MEM('o003464, 16'o104463);
`MEM('o003466, 16'o005201);
`MEM('o003470, 16'o010103);
`MEM('o003472, 16'o012701);
`MEM('o003474, 16'o013540);
`MEM('o003476, 16'o104472);
`MEM('o003500, 16'o104470);
`MEM('o003502, 16'o001402);
`MEM('o003504, 16'o005301);
`MEM('o003506, 16'o000652);
`MEM('o003510, 16'o104516);
`MEM('o003512, 16'o012701);
`MEM('o003514, 16'o013540);
`MEM('o003516, 16'o160103);
`MEM('o003520, 16'o010346);
`MEM('o003522, 16'o104410);
`MEM('o003524, 16'o005700);
`MEM('o003526, 16'o001436);
`MEM('o003530, 16'o020027);
`MEM('o003532, 16'o017777);
`MEM('o003534, 16'o003033);
`MEM('o003536, 16'o104474);
`MEM('o003540, 16'o001001);
`MEM('o003542, 16'o104476);
`MEM('o003544, 16'o012603);
`MEM('o003546, 16'o104516);
`MEM('o003550, 16'o010300);
`MEM('o003552, 16'o104504);
`MEM('o003554, 16'o103003);
`MEM('o003556, 16'o104401);
`MEM('o003560, 16'o060005);
`MEM('o003562, 16'o000410);
`MEM('o003564, 16'o020105);
`MEM('o003566, 16'o103374);
`MEM('o003570, 16'o010502);
`MEM('o003572, 16'o060005);
`MEM('o003574, 16'o010504);
`MEM('o003576, 16'o114244);
`MEM('o003600, 16'o020102);
`MEM('o003602, 16'o101775);
`MEM('o003604, 16'o012702);
`MEM('o003606, 16'o013540);
`MEM('o003610, 16'o111221);
`MEM('o003612, 16'o122227);
`MEM('o003614, 16'o000012);
`MEM('o003616, 16'o001374);
`MEM('o003620, 16'o000167);
`MEM('o003622, 16'o177160);
`MEM('o003624, 16'o104441);
`MEM('o003626, 16'o044514);
`MEM('o003630, 16'o052123);
`MEM('o003632, 16'o046044);
`MEM('o003634, 16'o052105);
`MEM('o003636, 16'o051044);
`MEM('o003640, 16'o040505);
`MEM('o003642, 16'o022104);
`MEM('o003644, 16'o042522);
`MEM('o003646, 16'o022115);
`MEM('o003650, 16'o052522);
`MEM('o003652, 16'o022116);
`MEM('o003654, 16'o042522);
`MEM('o003656, 16'o052123);
`MEM('o003660, 16'o051117);
`MEM('o003662, 16'o022105);
`MEM('o003664, 16'o042522);
`MEM('o003666, 16'o052524);
`MEM('o003670, 16'o047122);
`MEM('o003672, 16'o042044);
`MEM('o003674, 16'o052101);
`MEM('o003676, 16'o022101);
`MEM('o003700, 16'o044504);
`MEM('o003702, 16'o022115);
`MEM('o003704, 16'o042504);
`MEM('o003706, 16'o042514);
`MEM('o003710, 16'o042524);
`MEM('o003712, 16'o050044);
`MEM('o003714, 16'o044522);
`MEM('o003716, 16'o052116);
`MEM('o003720, 16'o043444);
`MEM('o003722, 16'o051517);
`MEM('o003724, 16'o041125);
`MEM('o003726, 16'o043444);
`MEM('o003730, 16'o052117);
`MEM('o003732, 16'o022117);
`MEM('o003734, 16'o043111);
`MEM('o003736, 16'o043044);
`MEM('o003740, 16'o051117);
`MEM('o003742, 16'o047044);
`MEM('o003744, 16'o054105);
`MEM('o003746, 16'o022124);
`MEM('o003750, 16'o047111);
`MEM('o003752, 16'o052520);
`MEM('o003754, 16'o022124);
`MEM('o003756, 16'o040523);
`MEM('o003760, 16'o042526);
`MEM('o003762, 16'o051444);
`MEM('o003764, 16'o047524);
`MEM('o003766, 16'o022120);
`MEM('o003770, 16'o047105);
`MEM('o003772, 16'o022104);
`MEM('o003774, 16'o042504);
`MEM('o003776, 16'o022106);
`MEM('o004000, 16'o046117);
`MEM('o004002, 16'o022104);
`MEM('o004004, 16'o040522);
`MEM('o004006, 16'o042116);
`MEM('o004010, 16'o046517);
`MEM('o004012, 16'o055111);
`MEM('o004014, 16'o022105);
`MEM('o004016, 16'o000044);
`MEM('o004020, 16'o002440);
`MEM('o004022, 16'o006070);
`MEM('o004024, 16'o007150);
`MEM('o004026, 16'o006324);
`MEM('o004030, 16'o004150);
`MEM('o004032, 16'o004240);
`MEM('o004034, 16'o004246);
`MEM('o004036, 16'o006324);
`MEM('o004040, 16'o004332);
`MEM('o004042, 16'o002670);
`MEM('o004044, 16'o006430);
`MEM('o004046, 16'o004204);
`MEM('o004050, 16'o004216);
`MEM('o004052, 16'o006140);
`MEM('o004054, 16'o007302);
`MEM('o004056, 16'o007620);
`MEM('o004060, 16'o006660);
`MEM('o004062, 16'o002060);
`MEM('o004064, 16'o004106);
`MEM('o004066, 16'o004106);
`MEM('o004070, 16'o004474);
`MEM('o004072, 16'o002072);
`MEM('o004074, 16'o010054);
`MEM('o004076, 16'o042522);
`MEM('o004100, 16'o042101);
`MEM('o004102, 16'o006531);
`MEM('o004104, 16'o000012);
`MEM('o004106, 16'o104402);
`MEM('o004110, 16'o012700);
`MEM('o004112, 16'o004132);
`MEM('o004114, 16'o104466);
`MEM('o004116, 16'o104404);
`MEM('o004120, 16'o104402);
`MEM('o004122, 16'o005067);
`MEM('o004124, 16'o007532);
`MEM('o004126, 16'o000167);
`MEM('o004130, 16'o176760);
`MEM('o004132, 16'o052123);
`MEM('o004134, 16'o050117);
`MEM('o004136, 16'o040440);
`MEM('o004140, 16'o020124);
`MEM('o004142, 16'o044514);
`MEM('o004144, 16'o042516);
`MEM('o004146, 16'o000040);
`MEM('o004150, 16'o104516);
`MEM('o004152, 16'o005067);
`MEM('o004154, 16'o007502);
`MEM('o004156, 16'o016701);
`MEM('o004160, 16'o007500);
`MEM('o004162, 16'o005201);
`MEM('o004164, 16'o012767);
`MEM('o004166, 16'o013507);
`MEM('o004170, 16'o003656);
`MEM('o004172, 16'o012767);
`MEM('o004174, 16'o000001);
`MEM('o004176, 16'o007464);
`MEM('o004200, 16'o000167);
`MEM('o004202, 16'o176600);
`MEM('o004204, 16'o016700);
`MEM('o004206, 16'o007450);
`MEM('o004210, 16'o052700);
`MEM('o004212, 16'o020000);
`MEM('o004214, 16'o104512);
`MEM('o004216, 16'o104410);
`MEM('o004220, 16'o104474);
`MEM('o004222, 16'o001005);
`MEM('o004224, 16'o012767);
`MEM('o004226, 16'o000001);
`MEM('o004230, 16'o007432);
`MEM('o004232, 16'o000167);
`MEM('o004234, 16'o176574);
`MEM('o004236, 16'o104405);
`MEM('o004240, 16'o005067);
`MEM('o004242, 16'o007424);
`MEM('o004244, 16'o000507);
`MEM('o004246, 16'o005046);
`MEM('o004250, 16'o012704);
`MEM('o004252, 16'o020000);
`MEM('o004254, 16'o104534);
`MEM('o004256, 16'o001424);
`MEM('o004260, 16'o012700);
`MEM('o004262, 16'o017777);
`MEM('o004264, 16'o104514);
`MEM('o004266, 16'o001403);
`MEM('o004270, 16'o010316);
`MEM('o004272, 16'o005723);
`MEM('o004274, 16'o000773);
`MEM('o004276, 16'o012603);
`MEM('o004300, 16'o001413);
`MEM('o004302, 16'o011300);
`MEM('o004304, 16'o040400);
`MEM('o004306, 16'o005200);
`MEM('o004310, 16'o012704);
`MEM('o004312, 16'o000002);
`MEM('o004314, 16'o104520);
`MEM('o004316, 16'o020027);
`MEM('o004320, 16'o000001);
`MEM('o004322, 16'o001677);
`MEM('o004324, 16'o104474);
`MEM('o004326, 16'o000736);
`MEM('o004330, 16'o104411);
`MEM('o004332, 16'o104544);
`MEM('o004334, 16'o102427);
`MEM('o004336, 16'o001055);
`MEM('o004340, 16'o010446);
`MEM('o004342, 16'o104472);
`MEM('o004344, 16'o020227);
`MEM('o004346, 16'o000050);
`MEM('o004350, 16'o001021);
`MEM('o004352, 16'o104410);
`MEM('o004354, 16'o104524);
`MEM('o004356, 16'o001016);
`MEM('o004360, 16'o010046);
`MEM('o004362, 16'o000316);
`MEM('o004364, 16'o104472);
`MEM('o004366, 16'o120227);
`MEM('o004370, 16'o000054);
`MEM('o004372, 16'o001005);
`MEM('o004374, 16'o104410);
`MEM('o004376, 16'o104524);
`MEM('o004400, 16'o001005);
`MEM('o004402, 16'o050016);
`MEM('o004404, 16'o104472);
`MEM('o004406, 16'o020227);
`MEM('o004410, 16'o000051);
`MEM('o004412, 16'o001401);
`MEM('o004414, 16'o104433);
`MEM('o004416, 16'o012602);
`MEM('o004420, 16'o012600);
`MEM('o004422, 16'o010146);
`MEM('o004424, 16'o104512);
`MEM('o004426, 16'o010200);
`MEM('o004430, 16'o104512);
`MEM('o004432, 16'o010201);
`MEM('o004434, 16'o000301);
`MEM('o004436, 16'o104522);
`MEM('o004440, 16'o102413);
`MEM('o004442, 16'o104504);
`MEM('o004444, 16'o103411);
`MEM('o004446, 16'o060005);
`MEM('o004450, 16'o012601);
`MEM('o004452, 16'o104472);
`MEM('o004454, 16'o020227);
`MEM('o004456, 16'o000054);
`MEM('o004460, 16'o001724);
`MEM('o004462, 16'o005301);
`MEM('o004464, 16'o000167);
`MEM('o004466, 16'o176272);
`MEM('o004470, 16'o104435);
`MEM('o004472, 16'o104443);
`MEM('o004474, 16'o104540);
`MEM('o004476, 16'o020427);
`MEM('o004500, 16'o043116);
`MEM('o004502, 16'o001033);
`MEM('o004504, 16'o104472);
`MEM('o004506, 16'o104470);
`MEM('o004510, 16'o001430);
`MEM('o004512, 16'o102427);
`MEM('o004514, 16'o052702);
`MEM('o004516, 16'o060000);
`MEM('o004520, 16'o010200);
`MEM('o004522, 16'o104512);
`MEM('o004524, 16'o104472);
`MEM('o004526, 16'o020227);
`MEM('o004530, 16'o000050);
`MEM('o004532, 16'o001017);
`MEM('o004534, 16'o104526);
`MEM('o004536, 16'o102415);
`MEM('o004540, 16'o010400);
`MEM('o004542, 16'o104512);
`MEM('o004544, 16'o020227);
`MEM('o004546, 16'o000051);
`MEM('o004550, 16'o001010);
`MEM('o004552, 16'o104472);
`MEM('o004554, 16'o020227);
`MEM('o004556, 16'o000075);
`MEM('o004560, 16'o001004);
`MEM('o004562, 16'o010100);
`MEM('o004564, 16'o104512);
`MEM('o004566, 16'o104510);
`MEM('o004570, 16'o000735);
`MEM('o004572, 16'o104437);
`MEM('o004574, 16'o005000);
`MEM('o004576, 16'o104512);
`MEM('o004600, 16'o012746);
`MEM('o004602, 16'o177777);
`MEM('o004604, 16'o104504);
`MEM('o004606, 16'o103561);
`MEM('o004610, 16'o104472);
`MEM('o004612, 16'o020227);
`MEM('o004614, 16'o000053);
`MEM('o004616, 16'o001410);
`MEM('o004620, 16'o020227);
`MEM('o004622, 16'o000055);
`MEM('o004624, 16'o001006);
`MEM('o004626, 16'o010200);
`MEM('o004630, 16'o005002);
`MEM('o004632, 16'o005003);
`MEM('o004634, 16'o005004);
`MEM('o004636, 16'o000410);
`MEM('o004640, 16'o104472);
`MEM('o004642, 16'o020227);
`MEM('o004644, 16'o000050);
`MEM('o004646, 16'o001007);
`MEM('o004650, 16'o005046);
`MEM('o004652, 16'o005265);
`MEM('o004654, 16'o177776);
`MEM('o004656, 16'o000752);
`MEM('o004660, 16'o104542);
`MEM('o004662, 16'o010046);
`MEM('o004664, 16'o000765);
`MEM('o004666, 16'o005301);
`MEM('o004670, 16'o014546);
`MEM('o004672, 16'o004767);
`MEM('o004674, 16'o000302);
`MEM('o004676, 16'o012625);
`MEM('o004700, 16'o010246);
`MEM('o004702, 16'o104472);
`MEM('o004704, 16'o012700);
`MEM('o004706, 16'o005163);
`MEM('o004710, 16'o124002);
`MEM('o004712, 16'o001407);
`MEM('o004714, 16'o020027);
`MEM('o004716, 16'o005155);
`MEM('o004720, 16'o101373);
`MEM('o004722, 16'o005000);
`MEM('o004724, 16'o005301);
`MEM('o004726, 16'o012602);
`MEM('o004730, 16'o000402);
`MEM('o004732, 16'o010200);
`MEM('o004734, 16'o000774);
`MEM('o004736, 16'o005716);
`MEM('o004740, 16'o003457);
`MEM('o004742, 16'o010146);
`MEM('o004744, 16'o012701);
`MEM('o004746, 16'o005163);
`MEM('o004750, 16'o124100);
`MEM('o004752, 16'o001376);
`MEM('o004754, 16'o006201);
`MEM('o004756, 16'o010125);
`MEM('o004760, 16'o012701);
`MEM('o004762, 16'o005163);
`MEM('o004764, 16'o124166);
`MEM('o004766, 16'o000002);
`MEM('o004770, 16'o001375);
`MEM('o004772, 16'o006201);
`MEM('o004774, 16'o010125);
`MEM('o004776, 16'o012601);
`MEM('o005000, 16'o024545);
`MEM('o005002, 16'o002726);
`MEM('o005004, 16'o010025);
`MEM('o005006, 16'o012700);
`MEM('o005010, 16'o005163);
`MEM('o005012, 16'o124016);
`MEM('o005014, 16'o001376);
`MEM('o005016, 16'o162700);
`MEM('o005020, 16'o005156);
`MEM('o005022, 16'o006300);
`MEM('o005024, 16'o062700);
`MEM('o005026, 16'o005164);
`MEM('o005030, 16'o010025);
`MEM('o005032, 16'o005726);
`MEM('o005034, 16'o010600);
`MEM('o005036, 16'o104542);
`MEM('o005040, 16'o010146);
`MEM('o005042, 16'o010601);
`MEM('o005044, 16'o005721);
`MEM('o005046, 16'o014502);
`MEM('o005050, 16'o014546);
`MEM('o005052, 16'o004772);
`MEM('o005054, 16'o000000);
`MEM('o005056, 16'o012600);
`MEM('o005060, 16'o012601);
`MEM('o005062, 16'o062706);
`MEM('o005064, 16'o000006);
`MEM('o005066, 16'o012602);
`MEM('o005070, 16'o012603);
`MEM('o005072, 16'o012604);
`MEM('o005074, 16'o005716);
`MEM('o005076, 16'o003321);
`MEM('o005100, 16'o020027);
`MEM('o005102, 16'o000051);
`MEM('o005104, 16'o001410);
`MEM('o005106, 16'o005700);
`MEM('o005110, 16'o003263);
`MEM('o005112, 16'o005745);
`MEM('o005114, 16'o001003);
`MEM('o005116, 16'o005726);
`MEM('o005120, 16'o000257);
`MEM('o005122, 16'o000207);
`MEM('o005124, 16'o104417);
`MEM('o005126, 16'o005745);
`MEM('o005130, 16'o001003);
`MEM('o005132, 16'o005726);
`MEM('o005134, 16'o000262);
`MEM('o005136, 16'o000207);
`MEM('o005140, 16'o005716);
`MEM('o005142, 16'o002773);
`MEM('o005144, 16'o005726);
`MEM('o005146, 16'o005325);
`MEM('o005150, 16'o000653);
`MEM('o005152, 16'o104401);
`MEM('o005154, 16'o024400);
`MEM('o005156, 16'o026453);
`MEM('o005160, 16'o027452);
`MEM('o005162, 16'o000136);
`MEM('o005164, 16'o012216);
`MEM('o005166, 16'o012442);
`MEM('o005170, 16'o012776);
`MEM('o005172, 16'o012550);
`MEM('o005174, 16'o013714);
`MEM('o005176, 16'o104467);
`MEM('o005200, 16'o010146);
`MEM('o005202, 16'o104472);
`MEM('o005204, 16'o104470);
`MEM('o005206, 16'o102417);
`MEM('o005210, 16'o001022);
`MEM('o005212, 16'o012601);
`MEM('o005214, 16'o162706);
`MEM('o005216, 16'o000006);
`MEM('o005220, 16'o010600);
`MEM('o005222, 16'o104406);
`MEM('o005224, 16'o102764);
`MEM('o005226, 16'o012602);
`MEM('o005230, 16'o012603);
`MEM('o005232, 16'o012604);
`MEM('o005234, 16'o000207);
`MEM('o005236, 16'o012002);
`MEM('o005240, 16'o012003);
`MEM('o005242, 16'o012004);
`MEM('o005244, 16'o000207);
`MEM('o005246, 16'o020227);
`MEM('o005250, 16'o000056);
`MEM('o005252, 16'o001757);
`MEM('o005254, 16'o000471);
`MEM('o005256, 16'o020227);
`MEM('o005260, 16'o000106);
`MEM('o005262, 16'o001473);
`MEM('o005264, 16'o012746);
`MEM('o005266, 16'o177700);
`MEM('o005270, 16'o041602);
`MEM('o005272, 16'o010200);
`MEM('o005274, 16'o104530);
`MEM('o005276, 16'o104530);
`MEM('o005300, 16'o104472);
`MEM('o005302, 16'o104470);
`MEM('o005304, 16'o102454);
`MEM('o005306, 16'o001453);
`MEM('o005310, 16'o041602);
`MEM('o005312, 16'o060200);
`MEM('o005314, 16'o104530);
`MEM('o005316, 16'o104530);
`MEM('o005320, 16'o104472);
`MEM('o005322, 16'o104470);
`MEM('o005324, 16'o102444);
`MEM('o005326, 16'o001443);
`MEM('o005330, 16'o042602);
`MEM('o005332, 16'o060200);
`MEM('o005334, 16'o012703);
`MEM('o005336, 16'o005734);
`MEM('o005340, 16'o022300);
`MEM('o005342, 16'o001404);
`MEM('o005344, 16'o020327);
`MEM('o005346, 16'o005762);
`MEM('o005350, 16'o103773);
`MEM('o005352, 16'o000552);
`MEM('o005354, 16'o104472);
`MEM('o005356, 16'o020227);
`MEM('o005360, 16'o000050);
`MEM('o005362, 16'o001146);
`MEM('o005364, 16'o016346);
`MEM('o005366, 16'o000024);
`MEM('o005370, 16'o104536);
`MEM('o005372, 16'o102023);
`MEM('o005374, 16'o012600);
`MEM('o005376, 16'o104542);
`MEM('o005400, 16'o010002);
`MEM('o005402, 16'o010600);
`MEM('o005404, 16'o010146);
`MEM('o005406, 16'o010001);
`MEM('o005410, 16'o162706);
`MEM('o005412, 16'o000006);
`MEM('o005414, 16'o010600);
`MEM('o005416, 16'o004712);
`MEM('o005420, 16'o012602);
`MEM('o005422, 16'o012603);
`MEM('o005424, 16'o012604);
`MEM('o005426, 16'o012601);
`MEM('o005430, 16'o062706);
`MEM('o005432, 16'o000010);
`MEM('o005434, 16'o000207);
`MEM('o005436, 16'o005726);
`MEM('o005440, 16'o000517);
`MEM('o005442, 16'o021627);
`MEM('o005444, 16'o017204);
`MEM('o005446, 16'o001036);
`MEM('o005450, 16'o000751);
`MEM('o005452, 16'o104472);
`MEM('o005454, 16'o020227);
`MEM('o005456, 16'o000116);
`MEM('o005460, 16'o001107);
`MEM('o005462, 16'o104472);
`MEM('o005464, 16'o104470);
`MEM('o005466, 16'o102504);
`MEM('o005470, 16'o001503);
`MEM('o005472, 16'o104534);
`MEM('o005474, 16'o001507);
`MEM('o005476, 16'o005000);
`MEM('o005500, 16'o052702);
`MEM('o005502, 16'o060000);
`MEM('o005504, 16'o010204);
`MEM('o005506, 16'o104514);
`MEM('o005510, 16'o001473);
`MEM('o005512, 16'o005723);
`MEM('o005514, 16'o012304);
`MEM('o005516, 16'o012346);
`MEM('o005520, 16'o104534);
`MEM('o005522, 16'o104514);
`MEM('o005524, 16'o001027);
`MEM('o005526, 16'o104472);
`MEM('o005530, 16'o020227);
`MEM('o005532, 16'o000050);
`MEM('o005534, 16'o001340);
`MEM('o005536, 16'o010446);
`MEM('o005540, 16'o104536);
`MEM('o005542, 16'o102401);
`MEM('o005544, 16'o104417);
`MEM('o005546, 16'o012600);
`MEM('o005550, 16'o010546);
`MEM('o005552, 16'o104512);
`MEM('o005554, 16'o005000);
`MEM('o005556, 16'o104512);
`MEM('o005560, 16'o104550);
`MEM('o005562, 16'o010146);
`MEM('o005564, 16'o016601);
`MEM('o005566, 16'o000004);
`MEM('o005570, 16'o104536);
`MEM('o005572, 16'o102764);
`MEM('o005574, 16'o012601);
`MEM('o005576, 16'o012605);
`MEM('o005600, 16'o022626);
`MEM('o005602, 16'o000207);
`MEM('o005604, 16'o022323);
`MEM('o005606, 16'o012600);
`MEM('o005610, 16'o012346);
`MEM('o005612, 16'o012346);
`MEM('o005614, 16'o012346);
`MEM('o005616, 16'o010346);
`MEM('o005620, 16'o010046);
`MEM('o005622, 16'o104472);
`MEM('o005624, 16'o020227);
`MEM('o005626, 16'o000050);
`MEM('o005630, 16'o001036);
`MEM('o005632, 16'o104536);
`MEM('o005634, 16'o102343);
`MEM('o005636, 16'o010100);
`MEM('o005640, 16'o016601);
`MEM('o005642, 16'o000002);
`MEM('o005644, 16'o010441);
`MEM('o005646, 16'o010341);
`MEM('o005650, 16'o010241);
`MEM('o005652, 16'o012601);
`MEM('o005654, 16'o010046);
`MEM('o005656, 16'o104536);
`MEM('o005660, 16'o102731);
`MEM('o005662, 16'o012601);
`MEM('o005664, 16'o012600);
`MEM('o005666, 16'o012640);
`MEM('o005670, 16'o012640);
`MEM('o005672, 16'o012640);
`MEM('o005674, 16'o005726);
`MEM('o005676, 16'o000207);
`MEM('o005700, 16'o012601);
`MEM('o005702, 16'o104544);
`MEM('o005704, 16'o102403);
`MEM('o005706, 16'o001402);
`MEM('o005710, 16'o000167);
`MEM('o005712, 16'o177322);
`MEM('o005714, 16'o104767);
`MEM('o005716, 16'o005002);
`MEM('o005720, 16'o005003);
`MEM('o005722, 16'o005004);
`MEM('o005724, 16'o000207);
`MEM('o005726, 16'o062706);
`MEM('o005730, 16'o000012);
`MEM('o005732, 16'o000762);
`MEM('o005734, 16'o060602);
`MEM('o005736, 16'o010537);
`MEM('o005740, 16'o003756);
`MEM('o005742, 16'o016300);
`MEM('o005744, 16'o037343);
`MEM('o005746, 16'o002553);
`MEM('o005750, 16'o061246);
`MEM('o005752, 16'o027634);
`MEM('o005754, 16'o056434);
`MEM('o005756, 16'o060472);
`MEM('o005760, 16'o016266);
`MEM('o005762, 16'o015020);
`MEM('o005764, 16'o015162);
`MEM('o005766, 16'o015260);
`MEM('o005770, 16'o014260);
`MEM('o005772, 16'o013764);
`MEM('o005774, 16'o012470);
`MEM('o005776, 16'o015642);
`MEM('o006000, 16'o013372);
`MEM('o006002, 16'o010004);
`MEM('o006004, 16'o012522);
`MEM('o006006, 16'o017204);
`MEM('o006010, 16'o104526);
`MEM('o006012, 16'o102422);
`MEM('o006014, 16'o005301);
`MEM('o006016, 16'o005000);
`MEM('o006020, 16'o104534);
`MEM('o006022, 16'o001415);
`MEM('o006024, 16'o104514);
`MEM('o006026, 16'o001413);
`MEM('o006030, 16'o021627);
`MEM('o006032, 16'o004334);
`MEM('o006034, 16'o001413);
`MEM('o006036, 16'o005723);
`MEM('o006040, 16'o121127);
`MEM('o006042, 16'o000050);
`MEM('o006044, 16'o001006);
`MEM('o006046, 16'o005201);
`MEM('o006050, 16'o010446);
`MEM('o006052, 16'o104532);
`MEM('o006054, 16'o012604);
`MEM('o006056, 16'o005700);
`MEM('o006060, 16'o000207);
`MEM('o006062, 16'o005723);
`MEM('o006064, 16'o010300);
`MEM('o006066, 16'o000207);
`MEM('o006070, 16'o104544);
`MEM('o006072, 16'o102420);
`MEM('o006074, 16'o001002);
`MEM('o006076, 16'o010400);
`MEM('o006100, 16'o104546);
`MEM('o006102, 16'o010046);
`MEM('o006104, 16'o104472);
`MEM('o006106, 16'o020227);
`MEM('o006110, 16'o000075);
`MEM('o006112, 16'o001010);
`MEM('o006114, 16'o104536);
`MEM('o006116, 16'o102407);
`MEM('o006120, 16'o012600);
`MEM('o006122, 16'o010220);
`MEM('o006124, 16'o010320);
`MEM('o006126, 16'o010420);
`MEM('o006130, 16'o000167);
`MEM('o006132, 16'o174626);
`MEM('o006134, 16'o104421);
`MEM('o006136, 16'o104417);
`MEM('o006140, 16'o104536);
`MEM('o006142, 16'o102775);
`MEM('o006144, 16'o104542);
`MEM('o006146, 16'o104540);
`MEM('o006150, 16'o020227);
`MEM('o006152, 16'o000076);
`MEM('o006154, 16'o001405);
`MEM('o006156, 16'o020227);
`MEM('o006160, 16'o000075);
`MEM('o006162, 16'o001402);
`MEM('o006164, 16'o005301);
`MEM('o006166, 16'o105004);
`MEM('o006170, 16'o012702);
`MEM('o006172, 16'o006250);
`MEM('o006174, 16'o020422);
`MEM('o006176, 16'o001404);
`MEM('o006200, 16'o020227);
`MEM('o006202, 16'o006264);
`MEM('o006204, 16'o103773);
`MEM('o006206, 16'o104423);
`MEM('o006210, 16'o062702);
`MEM('o006212, 16'o171526);
`MEM('o006214, 16'o006302);
`MEM('o006216, 16'o062702);
`MEM('o006220, 16'o006264);
`MEM('o006222, 16'o010246);
`MEM('o006224, 16'o104536);
`MEM('o006226, 16'o102743);
`MEM('o006230, 16'o010146);
`MEM('o006232, 16'o010601);
`MEM('o006234, 16'o022121);
`MEM('o006236, 16'o104542);
`MEM('o006240, 16'o010600);
`MEM('o006242, 16'o104434);
`MEM('o006244, 16'o000176);
`MEM('o006246, 16'o000010);
`MEM('o006250, 16'o036076);
`MEM('o006252, 16'o036075);
`MEM('o006254, 16'o036000);
`MEM('o006256, 16'o037075);
`MEM('o006260, 16'o037000);
`MEM('o006262, 16'o036400);
`MEM('o006264, 16'o001023);
`MEM('o006266, 16'o000411);
`MEM('o006270, 16'o003421);
`MEM('o006272, 16'o000407);
`MEM('o006274, 16'o002417);
`MEM('o006276, 16'o000405);
`MEM('o006300, 16'o002015);
`MEM('o006302, 16'o000403);
`MEM('o006304, 16'o003013);
`MEM('o006306, 16'o000401);
`MEM('o006310, 16'o001411);
`MEM('o006312, 16'o062706);
`MEM('o006314, 16'o000006);
`MEM('o006316, 16'o012601);
`MEM('o006320, 16'o062706);
`MEM('o006322, 16'o000010);
`MEM('o006324, 16'o104502);
`MEM('o006326, 16'o005301);
`MEM('o006330, 16'o000167);
`MEM('o006332, 16'o174426);
`MEM('o006334, 16'o062706);
`MEM('o006336, 16'o000006);
`MEM('o006340, 16'o012601);
`MEM('o006342, 16'o062706);
`MEM('o006344, 16'o000010);
`MEM('o006346, 16'o104540);
`MEM('o006350, 16'o020427);
`MEM('o006352, 16'o052110);
`MEM('o006354, 16'o001015);
`MEM('o006356, 16'o104540);
`MEM('o006360, 16'o020427);
`MEM('o006362, 16'o042516);
`MEM('o006364, 16'o001020);
`MEM('o006366, 16'o104472);
`MEM('o006370, 16'o005301);
`MEM('o006372, 16'o104470);
`MEM('o006374, 16'o102403);
`MEM('o006376, 16'o001013);
`MEM('o006400, 16'o000167);
`MEM('o006402, 16'o175612);
`MEM('o006404, 16'o000167);
`MEM('o006406, 16'o174624);
`MEM('o006410, 16'o020427);
`MEM('o006412, 16'o043517);
`MEM('o006414, 16'o001004);
`MEM('o006416, 16'o104540);
`MEM('o006420, 16'o020427);
`MEM('o006422, 16'o052117);
`MEM('o006424, 16'o001765);
`MEM('o006426, 16'o104425);
`MEM('o006430, 16'o005046);
`MEM('o006432, 16'o012700);
`MEM('o006434, 16'o000034);
`MEM('o006436, 16'o104504);
`MEM('o006440, 16'o103506);
`MEM('o006442, 16'o104472);
`MEM('o006444, 16'o120227);
`MEM('o006446, 16'o000054);
`MEM('o006450, 16'o001434);
`MEM('o006452, 16'o120227);
`MEM('o006454, 16'o000073);
`MEM('o006456, 16'o001452);
`MEM('o006460, 16'o120227);
`MEM('o006462, 16'o000042);
`MEM('o006464, 16'o001453);
`MEM('o006466, 16'o120227);
`MEM('o006470, 16'o000072);
`MEM('o006472, 16'o001463);
`MEM('o006474, 16'o120227);
`MEM('o006476, 16'o000012);
`MEM('o006500, 16'o001460);
`MEM('o006502, 16'o005716);
`MEM('o006504, 16'o002442);
`MEM('o006506, 16'o005301);
`MEM('o006510, 16'o104536);
`MEM('o006512, 16'o102437);
`MEM('o006514, 16'o010146);
`MEM('o006516, 16'o004767);
`MEM('o006520, 16'o002174);
`MEM('o006522, 16'o010600);
`MEM('o006524, 16'o104466);
`MEM('o006526, 16'o062706);
`MEM('o006530, 16'o000024);
`MEM('o006532, 16'o012601);
`MEM('o006534, 16'o012716);
`MEM('o006536, 16'o177777);
`MEM('o006540, 16'o000734);
`MEM('o006542, 16'o016700);
`MEM('o006544, 16'o005124);
`MEM('o006546, 16'o020027);
`MEM('o006550, 16'o000070);
`MEM('o006552, 16'o002402);
`MEM('o006554, 16'o104402);
`MEM('o006556, 16'o000412);
`MEM('o006560, 16'o005400);
`MEM('o006562, 16'o003003);
`MEM('o006564, 16'o062700);
`MEM('o006566, 16'o000016);
`MEM('o006570, 16'o000774);
`MEM('o006572, 16'o112702);
`MEM('o006574, 16'o000040);
`MEM('o006576, 16'o104400);
`MEM('o006600, 16'o005300);
`MEM('o006602, 16'o003375);
`MEM('o006604, 16'o012716);
`MEM('o006606, 16'o000001);
`MEM('o006610, 16'o000710);
`MEM('o006612, 16'o104427);
`MEM('o006614, 16'o112102);
`MEM('o006616, 16'o104400);
`MEM('o006620, 16'o121127);
`MEM('o006622, 16'o000012);
`MEM('o006624, 16'o001772);
`MEM('o006626, 16'o121127);
`MEM('o006630, 16'o000042);
`MEM('o006632, 16'o001370);
`MEM('o006634, 16'o005201);
`MEM('o006636, 16'o005016);
`MEM('o006640, 16'o000674);
`MEM('o006642, 16'o005726);
`MEM('o006644, 16'o003001);
`MEM('o006646, 16'o104402);
`MEM('o006650, 16'o005301);
`MEM('o006652, 16'o000167);
`MEM('o006654, 16'o174104);
`MEM('o006656, 16'o104401);
`MEM('o006660, 16'o005046);
`MEM('o006662, 16'o004767);
`MEM('o006664, 16'o000200);
`MEM('o006666, 16'o102001);
`MEM('o006670, 16'o104445);
`MEM('o006672, 16'o005046);
`MEM('o006674, 16'o010146);
`MEM('o006676, 16'o012702);
`MEM('o006700, 16'o000077);
`MEM('o006702, 16'o104400);
`MEM('o006704, 16'o104500);
`MEM('o006706, 16'o004767);
`MEM('o006710, 16'o000052);
`MEM('o006712, 16'o102422);
`MEM('o006714, 16'o003015);
`MEM('o006716, 16'o002416);
`MEM('o006720, 16'o012601);
`MEM('o006722, 16'o005726);
`MEM('o006724, 16'o005726);
`MEM('o006726, 16'o001376);
`MEM('o006730, 16'o005301);
`MEM('o006732, 16'o005767);
`MEM('o006734, 16'o004726);
`MEM('o006736, 16'o001002);
`MEM('o006740, 16'o112711);
`MEM('o006742, 16'o000012);
`MEM('o006744, 16'o000167);
`MEM('o006746, 16'o174012);
`MEM('o006750, 16'o104765);
`MEM('o006752, 16'o000751);
`MEM('o006754, 16'o104763);
`MEM('o006756, 16'o000747);
`MEM('o006760, 16'o104761);
`MEM('o006762, 16'o000745);
`MEM('o006764, 16'o010604);
`MEM('o006766, 16'o022424);
`MEM('o006770, 16'o005724);
`MEM('o006772, 16'o005724);
`MEM('o006774, 16'o001376);
`MEM('o006776, 16'o005744);
`MEM('o007000, 16'o014400);
`MEM('o007002, 16'o001425);
`MEM('o007004, 16'o010446);
`MEM('o007006, 16'o104406);
`MEM('o007010, 16'o102424);
`MEM('o007012, 16'o012604);
`MEM('o007014, 16'o121127);
`MEM('o007016, 16'o000054);
`MEM('o007020, 16'o001410);
`MEM('o007022, 16'o121127);
`MEM('o007024, 16'o000072);
`MEM('o007026, 16'o001407);
`MEM('o007030, 16'o121127);
`MEM('o007032, 16'o000012);
`MEM('o007034, 16'o001404);
`MEM('o007036, 16'o000262);
`MEM('o007040, 16'o000207);
`MEM('o007042, 16'o005201);
`MEM('o007044, 16'o000755);
`MEM('o007046, 16'o014400);
`MEM('o007050, 16'o001773);
`MEM('o007052, 16'o000270);
`MEM('o007054, 16'o000207);
`MEM('o007056, 16'o000257);
`MEM('o007060, 16'o000207);
`MEM('o007062, 16'o005726);
`MEM('o007064, 16'o000764);
`MEM('o007066, 16'o104544);
`MEM('o007070, 16'o102424);
`MEM('o007072, 16'o001002);
`MEM('o007074, 16'o010400);
`MEM('o007076, 16'o104546);
`MEM('o007100, 16'o012602);
`MEM('o007102, 16'o010046);
`MEM('o007104, 16'o012700);
`MEM('o007106, 16'o000004);
`MEM('o007110, 16'o104504);
`MEM('o007112, 16'o103415);
`MEM('o007114, 16'o010246);
`MEM('o007116, 16'o104472);
`MEM('o007120, 16'o120227);
`MEM('o007122, 16'o000054);
`MEM('o007124, 16'o001760);
`MEM('o007126, 16'o120227);
`MEM('o007130, 16'o000072);
`MEM('o007132, 16'o001404);
`MEM('o007134, 16'o120227);
`MEM('o007136, 16'o000012);
`MEM('o007140, 16'o001401);
`MEM('o007142, 16'o000262);
`MEM('o007144, 16'o000207);
`MEM('o007146, 16'o104401);
`MEM('o007150, 16'o012746);
`MEM('o007152, 16'o000001);
`MEM('o007154, 16'o005046);
`MEM('o007156, 16'o004767);
`MEM('o007160, 16'o177704);
`MEM('o007162, 16'o102001);
`MEM('o007164, 16'o104447);
`MEM('o007166, 16'o005046);
`MEM('o007170, 16'o010146);
`MEM('o007172, 16'o016701);
`MEM('o007174, 16'o004472);
`MEM('o007176, 16'o001003);
`MEM('o007200, 16'o016701);
`MEM('o007202, 16'o004456);
`MEM('o007204, 16'o000426);
`MEM('o007206, 16'o121127);
`MEM('o007210, 16'o000012);
`MEM('o007212, 16'o001423);
`MEM('o007214, 16'o004767);
`MEM('o007216, 16'o177544);
`MEM('o007220, 16'o102427);
`MEM('o007222, 16'o002413);
`MEM('o007224, 16'o010167);
`MEM('o007226, 16'o004440);
`MEM('o007230, 16'o012601);
`MEM('o007232, 16'o005726);
`MEM('o007234, 16'o005726);
`MEM('o007236, 16'o001376);
`MEM('o007240, 16'o005726);
`MEM('o007242, 16'o001776);
`MEM('o007244, 16'o005301);
`MEM('o007246, 16'o000167);
`MEM('o007250, 16'o173510);
`MEM('o007252, 16'o005724);
`MEM('o007254, 16'o005024);
`MEM('o007256, 16'o005714);
`MEM('o007260, 16'o001375);
`MEM('o007262, 16'o104534);
`MEM('o007264, 16'o122721);
`MEM('o007266, 16'o000147);
`MEM('o007270, 16'o001746);
`MEM('o007272, 16'o020103);
`MEM('o007274, 16'o103773);
`MEM('o007276, 16'o104451);
`MEM('o007300, 16'o104453);
`MEM('o007302, 16'o104526);
`MEM('o007304, 16'o020227);
`MEM('o007306, 16'o000075);
`MEM('o007310, 16'o001117);
`MEM('o007312, 16'o005000);
`MEM('o007314, 16'o010446);
`MEM('o007316, 16'o104534);
`MEM('o007320, 16'o104514);
`MEM('o007322, 16'o001003);
`MEM('o007324, 16'o010400);
`MEM('o007326, 16'o104546);
`MEM('o007330, 16'o000402);
`MEM('o007332, 16'o010300);
`MEM('o007334, 16'o022020);
`MEM('o007336, 16'o010046);
`MEM('o007340, 16'o005000);
`MEM('o007342, 16'o104534);
`MEM('o007344, 16'o052704);
`MEM('o007346, 16'o040000);
`MEM('o007350, 16'o104514);
`MEM('o007352, 16'o001407);
`MEM('o007354, 16'o010446);
`MEM('o007356, 16'o010146);
`MEM('o007360, 16'o012704);
`MEM('o007362, 16'o000020);
`MEM('o007364, 16'o104520);
`MEM('o007366, 16'o012601);
`MEM('o007370, 16'o012604);
`MEM('o007372, 16'o010400);
`MEM('o007374, 16'o104512);
`MEM('o007376, 16'o016700);
`MEM('o007400, 16'o004256);
`MEM('o007402, 16'o104512);
`MEM('o007404, 16'o104536);
`MEM('o007406, 16'o011600);
`MEM('o007410, 16'o010220);
`MEM('o007412, 16'o010320);
`MEM('o007414, 16'o010420);
`MEM('o007416, 16'o104540);
`MEM('o007420, 16'o020427);
`MEM('o007422, 16'o052117);
`MEM('o007424, 16'o001051);
`MEM('o007426, 16'o104536);
`MEM('o007430, 16'o104550);
`MEM('o007432, 16'o121127);
`MEM('o007434, 16'o000123);
`MEM('o007436, 16'o001013);
`MEM('o007440, 16'o104540);
`MEM('o007442, 16'o020427);
`MEM('o007444, 16'o051524);
`MEM('o007446, 16'o001040);
`MEM('o007450, 16'o104540);
`MEM('o007452, 16'o020427);
`MEM('o007454, 16'o042520);
`MEM('o007456, 16'o001034);
`MEM('o007460, 16'o104536);
`MEM('o007462, 16'o104550);
`MEM('o007464, 16'o000406);
`MEM('o007466, 16'o005002);
`MEM('o007470, 16'o012703);
`MEM('o007472, 16'o040000);
`MEM('o007474, 16'o012704);
`MEM('o007476, 16'o100001);
`MEM('o007500, 16'o000770);
`MEM('o007502, 16'o011600);
`MEM('o007504, 16'o010146);
`MEM('o007506, 16'o010501);
`MEM('o007510, 16'o162701);
`MEM('o007512, 16'o000014);
`MEM('o007514, 16'o010146);
`MEM('o007516, 16'o104434);
`MEM('o007520, 16'o001406);
`MEM('o007522, 16'o002413);
`MEM('o007524, 16'o012601);
`MEM('o007526, 16'o005761);
`MEM('o007530, 16'o000010);
`MEM('o007532, 16'o002413);
`MEM('o007534, 16'o000401);
`MEM('o007536, 16'o005726);
`MEM('o007540, 16'o012601);
`MEM('o007542, 16'o022626);
`MEM('o007544, 16'o000167);
`MEM('o007546, 16'o173212);
`MEM('o007550, 16'o104455);
`MEM('o007552, 16'o012601);
`MEM('o007554, 16'o005761);
`MEM('o007556, 16'o000010);
`MEM('o007560, 16'o002767);
`MEM('o007562, 16'o012601);
`MEM('o007564, 16'o005726);
`MEM('o007566, 16'o104534);
`MEM('o007570, 16'o122127);
`MEM('o007572, 16'o000157);
`MEM('o007574, 16'o001403);
`MEM('o007576, 16'o020103);
`MEM('o007600, 16'o103773);
`MEM('o007602, 16'o104457);
`MEM('o007604, 16'o104526);
`MEM('o007606, 16'o020416);
`MEM('o007610, 16'o001367);
`MEM('o007612, 16'o005726);
`MEM('o007614, 16'o005301);
`MEM('o007616, 16'o000752);
`MEM('o007620, 16'o005000);
`MEM('o007622, 16'o104526);
`MEM('o007624, 16'o010446);
`MEM('o007626, 16'o104534);
`MEM('o007630, 16'o104514);
`MEM('o007632, 16'o001451);
`MEM('o007634, 16'o010346);
`MEM('o007636, 16'o052704);
`MEM('o007640, 16'o040000);
`MEM('o007642, 16'o104534);
`MEM('o007644, 16'o104514);
`MEM('o007646, 16'o001443);
`MEM('o007650, 16'o010146);
`MEM('o007652, 16'o022323);
`MEM('o007654, 16'o010301);
`MEM('o007656, 16'o062701);
`MEM('o007660, 16'o000006);
`MEM('o007662, 16'o016600);
`MEM('o007664, 16'o000002);
`MEM('o007666, 16'o010346);
`MEM('o007670, 16'o022020);
`MEM('o007672, 16'o010046);
`MEM('o007674, 16'o104420);
`MEM('o007676, 16'o012600);
`MEM('o007700, 16'o011603);
`MEM('o007702, 16'o010301);
`MEM('o007704, 16'o005763);
`MEM('o007706, 16'o000010);
`MEM('o007710, 16'o100003);
`MEM('o007712, 16'o104434);
`MEM('o007714, 16'o003021);
`MEM('o007716, 16'o000402);
`MEM('o007720, 16'o104434);
`MEM('o007722, 16'o002416);
`MEM('o007724, 16'o012600);
`MEM('o007726, 16'o005726);
`MEM('o007730, 16'o010046);
`MEM('o007732, 16'o005740);
`MEM('o007734, 16'o011000);
`MEM('o007736, 16'o104474);
`MEM('o007740, 16'o104510);
`MEM('o007742, 16'o010104);
`MEM('o007744, 16'o012601);
`MEM('o007746, 16'o011600);
`MEM('o007750, 16'o010446);
`MEM('o007752, 16'o022020);
`MEM('o007754, 16'o000657);
`MEM('o007756, 16'o104461);
`MEM('o007760, 16'o012601);
`MEM('o007762, 16'o062701);
`MEM('o007764, 16'o000006);
`MEM('o007766, 16'o016600);
`MEM('o007770, 16'o000002);
`MEM('o007772, 16'o022020);
`MEM('o007774, 16'o104422);
`MEM('o007776, 16'o012601);
`MEM('o010000, 16'o022626);
`MEM('o010002, 16'o000704);
`MEM('o010004, 16'o010046);
`MEM('o010006, 16'o016700);
`MEM('o010010, 16'o000036);
`MEM('o010012, 16'o016701);
`MEM('o010014, 16'o000034);
`MEM('o010016, 16'o104416);
`MEM('o010020, 16'o042700);
`MEM('o010022, 16'o100000);
`MEM('o010024, 16'o010067);
`MEM('o010026, 16'o000020);
`MEM('o010030, 16'o010001);
`MEM('o010032, 16'o011600);
`MEM('o010034, 16'o104436);
`MEM('o010036, 16'o012600);
`MEM('o010040, 16'o162760);
`MEM('o010042, 16'o000017);
`MEM('o010044, 16'o000004);
`MEM('o010046, 16'o000207);
`MEM('o010050, 16'o013507);
`MEM('o010052, 16'o000403);
`MEM('o010054, 16'o016767);
`MEM('o010056, 16'o003630);
`MEM('o010060, 16'o177766);
`MEM('o010062, 16'o052767);
`MEM('o010064, 16'o000001);
`MEM('o010066, 16'o177760);
`MEM('o010070, 16'o000167);
`MEM('o010072, 16'o172666);
`MEM('o010074, 16'o010546);
`MEM('o010076, 16'o010046);
`MEM('o010100, 16'o005020);
`MEM('o010102, 16'o005020);
`MEM('o010104, 16'o005010);
`MEM('o010106, 16'o005046);
`MEM('o010110, 16'o005046);
`MEM('o010112, 16'o005046);
`MEM('o010114, 16'o104472);
`MEM('o010116, 16'o122702);
`MEM('o010120, 16'o000105);
`MEM('o010122, 16'o001474);
`MEM('o010124, 16'o122702);
`MEM('o010126, 16'o000055);
`MEM('o010130, 16'o001512);
`MEM('o010132, 16'o122702);
`MEM('o010134, 16'o000053);
`MEM('o010136, 16'o001504);
`MEM('o010140, 16'o122702);
`MEM('o010142, 16'o000056);
`MEM('o010144, 16'o001473);
`MEM('o010146, 16'o104470);
`MEM('o010150, 16'o001125);
`MEM('o010152, 16'o162702);
`MEM('o010154, 16'o000060);
`MEM('o010156, 16'o010146);
`MEM('o010160, 16'o032766);
`MEM('o010162, 16'o000004);
`MEM('o010164, 16'o000002);
`MEM('o010166, 16'o001033);
`MEM('o010170, 16'o162706);
`MEM('o010172, 16'o000006);
`MEM('o010174, 16'o010600);
`MEM('o010176, 16'o010201);
`MEM('o010200, 16'o104436);
`MEM('o010202, 16'o016600);
`MEM('o010204, 16'o000016);
`MEM('o010206, 16'o012701);
`MEM('o010210, 16'o010660);
`MEM('o010212, 16'o104430);
`MEM('o010214, 16'o102526);
`MEM('o010216, 16'o016600);
`MEM('o010220, 16'o000016);
`MEM('o010222, 16'o010601);
`MEM('o010224, 16'o104420);
`MEM('o010226, 16'o032766);
`MEM('o010230, 16'o000010);
`MEM('o010232, 16'o000010);
`MEM('o010234, 16'o001402);
`MEM('o010236, 16'o005366);
`MEM('o010240, 16'o000012);
`MEM('o010242, 16'o062706);
`MEM('o010244, 16'o000006);
`MEM('o010246, 16'o012601);
`MEM('o010250, 16'o052716);
`MEM('o010252, 16'o000001);
`MEM('o010254, 16'o000464);
`MEM('o010256, 16'o010246);
`MEM('o010260, 16'o016603);
`MEM('o010262, 16'o000010);
`MEM('o010264, 16'o012705);
`MEM('o010266, 16'o000012);
`MEM('o010270, 16'o005002);
`MEM('o010272, 16'o005004);
`MEM('o010274, 16'o020327);
`MEM('o010276, 16'o001724);
`MEM('o010300, 16'o003100);
`MEM('o010302, 16'o104462);
`MEM('o010304, 16'o062603);
`MEM('o010306, 16'o010366);
`MEM('o010310, 16'o000006);
`MEM('o010312, 16'o000755);
`MEM('o010314, 16'o032716);
`MEM('o010316, 16'o000004);
`MEM('o010320, 16'o001061);
`MEM('o010322, 16'o052716);
`MEM('o010324, 16'o000004);
`MEM('o010326, 16'o042716);
`MEM('o010330, 16'o000001);
`MEM('o010332, 16'o000435);
`MEM('o010334, 16'o032716);
`MEM('o010336, 16'o000014);
`MEM('o010340, 16'o001051);
`MEM('o010342, 16'o052716);
`MEM('o010344, 16'o000010);
`MEM('o010346, 16'o000427);
`MEM('o010350, 16'o042716);
`MEM('o010352, 16'o000400);
`MEM('o010354, 16'o000401);
`MEM('o010356, 16'o052716);
`MEM('o010360, 16'o000400);
`MEM('o010362, 16'o032716);
`MEM('o010364, 16'o000004);
`MEM('o010366, 16'o001020);
`MEM('o010370, 16'o032716);
`MEM('o010372, 16'o000001);
`MEM('o010374, 16'o001013);
`MEM('o010376, 16'o032716);
`MEM('o010400, 16'o000030);
`MEM('o010402, 16'o001030);
`MEM('o010404, 16'o052716);
`MEM('o010406, 16'o000020);
`MEM('o010410, 16'o032716);
`MEM('o010412, 16'o000400);
`MEM('o010414, 16'o001404);
`MEM('o010416, 16'o052716);
`MEM('o010420, 16'o000100);
`MEM('o010422, 16'o000401);
`MEM('o010424, 16'o000430);
`MEM('o010426, 16'o000632);
`MEM('o010430, 16'o032716);
`MEM('o010432, 16'o000001);
`MEM('o010434, 16'o001373);
`MEM('o010436, 16'o031627);
`MEM('o010440, 16'o000040);
`MEM('o010442, 16'o001010);
`MEM('o010444, 16'o052716);
`MEM('o010446, 16'o000040);
`MEM('o010450, 16'o032716);
`MEM('o010452, 16'o000400);
`MEM('o010454, 16'o001764);
`MEM('o010456, 16'o052716);
`MEM('o010460, 16'o000200);
`MEM('o010462, 16'o000761);
`MEM('o010464, 16'o052716);
`MEM('o010466, 16'o000002);
`MEM('o010470, 16'o000755);
`MEM('o010472, 16'o062706);
`MEM('o010474, 16'o000010);
`MEM('o010476, 16'o012601);
`MEM('o010500, 16'o000771);
`MEM('o010502, 16'o022626);
`MEM('o010504, 16'o000767);
`MEM('o010506, 16'o010146);
`MEM('o010510, 16'o032766);
`MEM('o010512, 16'o000100);
`MEM('o010514, 16'o000002);
`MEM('o010516, 16'o001404);
`MEM('o010520, 16'o016600);
`MEM('o010522, 16'o000010);
`MEM('o010524, 16'o010001);
`MEM('o010526, 16'o104424);
`MEM('o010530, 16'o032766);
`MEM('o010532, 16'o000200);
`MEM('o010534, 16'o000002);
`MEM('o010536, 16'o001407);
`MEM('o010540, 16'o005466);
`MEM('o010542, 16'o000006);
`MEM('o010544, 16'o102004);
`MEM('o010546, 16'o052766);
`MEM('o010550, 16'o000002);
`MEM('o010552, 16'o000002);
`MEM('o010554, 16'o000426);
`MEM('o010556, 16'o066666);
`MEM('o010560, 16'o000004);
`MEM('o010562, 16'o000006);
`MEM('o010564, 16'o001422);
`MEM('o010566, 16'o002411);
`MEM('o010570, 16'o016600);
`MEM('o010572, 16'o000010);
`MEM('o010574, 16'o012701);
`MEM('o010576, 16'o010660);
`MEM('o010600, 16'o104430);
`MEM('o010602, 16'o005366);
`MEM('o010604, 16'o000006);
`MEM('o010606, 16'o003370);
`MEM('o010610, 16'o000410);
`MEM('o010612, 16'o016600);
`MEM('o010614, 16'o000010);
`MEM('o010616, 16'o012701);
`MEM('o010620, 16'o010660);
`MEM('o010622, 16'o104426);
`MEM('o010624, 16'o005266);
`MEM('o010626, 16'o000006);
`MEM('o010630, 16'o002770);
`MEM('o010632, 16'o012601);
`MEM('o010634, 16'o005301);
`MEM('o010636, 16'o012604);
`MEM('o010640, 16'o062706);
`MEM('o010642, 16'o000006);
`MEM('o010644, 16'o012605);
`MEM('o010646, 16'o032704);
`MEM('o010650, 16'o000002);
`MEM('o010652, 16'o001401);
`MEM('o010654, 16'o000262);
`MEM('o010656, 16'o000207);
`MEM('o010660, 16'o000000);
`MEM('o010662, 16'o050000);
`MEM('o010664, 16'o100004);
`MEM('o010666, 16'o000000);
`MEM('o010670, 16'o040000);
`MEM('o010672, 16'o100001);
`MEM('o010674, 16'o000000);
`MEM('o010676, 16'o075022);
`MEM('o010700, 16'o100024);
`MEM('o010702, 16'o040000);
`MEM('o010704, 16'o046113);
`MEM('o010706, 16'o100030);
`MEM('o010710, 16'o000000);
`MEM('o010712, 16'o040000);
`MEM('o010714, 16'o100000);
`MEM('o010716, 16'o012700);
`MEM('o010720, 16'o000012);
`MEM('o010722, 16'o005046);
`MEM('o010724, 16'o005300);
`MEM('o010726, 16'o003375);
`MEM('o010730, 16'o104542);
`MEM('o010732, 16'o012766);
`MEM('o010734, 16'o030040);
`MEM('o010736, 16'o000010);
`MEM('o010740, 16'o112766);
`MEM('o010742, 16'o000040);
`MEM('o010744, 16'o000012);
`MEM('o010746, 16'o005703);
`MEM('o010750, 16'o001546);
`MEM('o010752, 16'o003006);
`MEM('o010754, 16'o010600);
`MEM('o010756, 16'o010001);
`MEM('o010760, 16'o104424);
`MEM('o010762, 16'o112766);
`MEM('o010764, 16'o000055);
`MEM('o010766, 16'o000010);
`MEM('o010770, 16'o012701);
`MEM('o010772, 16'o010674);
`MEM('o010774, 16'o010600);
`MEM('o010776, 16'o104434);
`MEM('o011000, 16'o003014);
`MEM('o011002, 16'o012700);
`MEM('o011004, 16'o010702);
`MEM('o011006, 16'o010601);
`MEM('o011010, 16'o104434);
`MEM('o011012, 16'o002416);
`MEM('o011014, 16'o012701);
`MEM('o011016, 16'o010660);
`MEM('o011020, 16'o010600);
`MEM('o011022, 16'o104426);
`MEM('o011024, 16'o005266);
`MEM('o011026, 16'o000006);
`MEM('o011030, 16'o000764);
`MEM('o011032, 16'o012701);
`MEM('o011034, 16'o010660);
`MEM('o011036, 16'o010600);
`MEM('o011040, 16'o104430);
`MEM('o011042, 16'o005366);
`MEM('o011044, 16'o000006);
`MEM('o011046, 16'o000750);
`MEM('o011050, 16'o012701);
`MEM('o011052, 16'o010710);
`MEM('o011054, 16'o010600);
`MEM('o011056, 16'o104420);
`MEM('o011060, 16'o162766);
`MEM('o011062, 16'o100037);
`MEM('o011064, 16'o000004);
`MEM('o011066, 16'o006266);
`MEM('o011070, 16'o000002);
`MEM('o011072, 16'o006016);
`MEM('o011074, 16'o005266);
`MEM('o011076, 16'o000004);
`MEM('o011100, 16'o001372);
`MEM('o011102, 16'o010600);
`MEM('o011104, 16'o062700);
`MEM('o011106, 16'o000016);
`MEM('o011110, 16'o010601);
`MEM('o011112, 16'o010046);
`MEM('o011114, 16'o104414);
`MEM('o011116, 16'o012600);
`MEM('o011120, 16'o062700);
`MEM('o011122, 16'o000003);
`MEM('o011124, 16'o122710);
`MEM('o011126, 16'o000040);
`MEM('o011130, 16'o001403);
`MEM('o011132, 16'o005266);
`MEM('o011134, 16'o000006);
`MEM('o011136, 16'o000401);
`MEM('o011140, 16'o005200);
`MEM('o011142, 16'o062766);
`MEM('o011144, 16'o000007);
`MEM('o011146, 16'o000006);
`MEM('o011150, 16'o012701);
`MEM('o011152, 16'o000010);
`MEM('o011154, 16'o010002);
`MEM('o011156, 16'o062702);
`MEM('o011160, 16'o000007);
`MEM('o011162, 16'o005301);
`MEM('o011164, 16'o122742);
`MEM('o011166, 16'o000060);
`MEM('o011170, 16'o001774);
`MEM('o011172, 16'o010604);
`MEM('o011174, 16'o062704);
`MEM('o011176, 16'o000011);
`MEM('o011200, 16'o022766);
`MEM('o011202, 16'o000010);
`MEM('o011204, 16'o000006);
`MEM('o011206, 16'o003450);
`MEM('o011210, 16'o022766);
`MEM('o011212, 16'o177770);
`MEM('o011214, 16'o000006);
`MEM('o011216, 16'o002044);
`MEM('o011220, 16'o010103);
`MEM('o011222, 16'o005403);
`MEM('o011224, 16'o066603);
`MEM('o011226, 16'o000006);
`MEM('o011230, 16'o062703);
`MEM('o011232, 16'o000007);
`MEM('o011234, 16'o002435);
`MEM('o011236, 16'o016603);
`MEM('o011240, 16'o000006);
`MEM('o011242, 16'o002415);
`MEM('o011244, 16'o003023);
`MEM('o011246, 16'o112724);
`MEM('o011250, 16'o000056);
`MEM('o011252, 16'o112024);
`MEM('o011254, 16'o020002);
`MEM('o011256, 16'o101775);
`MEM('o011260, 16'o112724);
`MEM('o011262, 16'o000040);
`MEM('o011264, 16'o105014);
`MEM('o011266, 16'o062706);
`MEM('o011270, 16'o000010);
`MEM('o011272, 16'o016607);
`MEM('o011274, 16'o000022);
`MEM('o011276, 16'o112724);
`MEM('o011300, 16'o000056);
`MEM('o011302, 16'o112724);
`MEM('o011304, 16'o000060);
`MEM('o011306, 16'o005203);
`MEM('o011310, 16'o002774);
`MEM('o011312, 16'o000757);
`MEM('o011314, 16'o112024);
`MEM('o011316, 16'o005303);
`MEM('o011320, 16'o003375);
`MEM('o011322, 16'o020002);
`MEM('o011324, 16'o101750);
`MEM('o011326, 16'o000754);
`MEM('o011330, 16'o112724);
`MEM('o011332, 16'o000056);
`MEM('o011334, 16'o112024);
`MEM('o011336, 16'o020002);
`MEM('o011340, 16'o101775);
`MEM('o011342, 16'o112724);
`MEM('o011344, 16'o000105);
`MEM('o011346, 16'o062706);
`MEM('o011350, 16'o000006);
`MEM('o011352, 16'o011601);
`MEM('o011354, 16'o010600);
`MEM('o011356, 16'o062700);
`MEM('o011360, 16'o000014);
`MEM('o011362, 16'o010046);
`MEM('o011364, 16'o010446);
`MEM('o011366, 16'o104412);
`MEM('o011370, 16'o012604);
`MEM('o011372, 16'o012600);
`MEM('o011374, 16'o122027);
`MEM('o011376, 16'o000040);
`MEM('o011400, 16'o001775);
`MEM('o011402, 16'o124027);
`MEM('o011404, 16'o000055);
`MEM('o011406, 16'o001402);
`MEM('o011410, 16'o112724);
`MEM('o011412, 16'o000040);
`MEM('o011414, 16'o112024);
`MEM('o011416, 16'o121027);
`MEM('o011420, 16'o000040);
`MEM('o011422, 16'o001374);
`MEM('o011424, 16'o112724);
`MEM('o011426, 16'o000040);
`MEM('o011430, 16'o105014);
`MEM('o011432, 16'o005726);
`MEM('o011434, 16'o016607);
`MEM('o011436, 16'o000022);
`MEM('o011440, 16'o005000);
`MEM('o011442, 16'o004767);
`MEM('o011444, 16'o167556);
`MEM('o011446, 16'o004767);
`MEM('o011450, 16'o166756);
`MEM('o011452, 16'o001013);
`MEM('o011454, 16'o162702);
`MEM('o011456, 16'o000060);
`MEM('o011460, 16'o006300);
`MEM('o011462, 16'o060002);
`MEM('o011464, 16'o006300);
`MEM('o011466, 16'o006300);
`MEM('o011470, 16'o060200);
`MEM('o011472, 16'o032700);
`MEM('o011474, 16'o160000);
`MEM('o011476, 16'o001761);
`MEM('o011500, 16'o104441);
`MEM('o011502, 16'o005301);
`MEM('o011504, 16'o000207);
`MEM('o011506, 16'o010046);
`MEM('o011510, 16'o005046);
`MEM('o011512, 16'o010146);
`MEM('o011514, 16'o002002);
`MEM('o011516, 16'o005166);
`MEM('o011520, 16'o000002);
`MEM('o011522, 16'o010601);
`MEM('o011524, 16'o162706);
`MEM('o011526, 16'o000014);
`MEM('o011530, 16'o010600);
`MEM('o011532, 16'o104414);
`MEM('o011534, 16'o010601);
`MEM('o011536, 16'o016600);
`MEM('o011540, 16'o000020);
`MEM('o011542, 16'o062701);
`MEM('o011544, 16'o000005);
`MEM('o011546, 16'o012702);
`MEM('o011550, 16'o000007);
`MEM('o011552, 16'o112120);
`MEM('o011554, 16'o005302);
`MEM('o011556, 16'o003375);
`MEM('o011560, 16'o062706);
`MEM('o011562, 16'o000022);
`MEM('o011564, 16'o000207);
`MEM('o011566, 16'o010546);
`MEM('o011570, 16'o010046);
`MEM('o011572, 16'o005046);
`MEM('o011574, 16'o012103);
`MEM('o011576, 16'o011102);
`MEM('o011600, 16'o002004);
`MEM('o011602, 16'o005402);
`MEM('o011604, 16'o005403);
`MEM('o011606, 16'o005602);
`MEM('o011610, 16'o005216);
`MEM('o011612, 16'o012705);
`MEM('o011614, 16'o000012);
`MEM('o011616, 16'o005004);
`MEM('o011620, 16'o012746);
`MEM('o011622, 16'o177777);
`MEM('o011624, 16'o005000);
`MEM('o011626, 16'o005001);
`MEM('o011630, 16'o104464);
`MEM('o011632, 16'o010146);
`MEM('o011634, 16'o050200);
`MEM('o011636, 16'o050300);
`MEM('o011640, 16'o005700);
`MEM('o011642, 16'o001370);
`MEM('o011644, 16'o010605);
`MEM('o011646, 16'o005204);
`MEM('o011650, 16'o005725);
`MEM('o011652, 16'o002375);
`MEM('o011654, 16'o005304);
`MEM('o011656, 16'o012703);
`MEM('o011660, 16'o000013);
`MEM('o011662, 16'o160403);
`MEM('o011664, 16'o005303);
`MEM('o011666, 16'o016500);
`MEM('o011670, 16'o000002);
`MEM('o011672, 16'o005703);
`MEM('o011674, 16'o003404);
`MEM('o011676, 16'o112720);
`MEM('o011700, 16'o000040);
`MEM('o011702, 16'o005303);
`MEM('o011704, 16'o000772);
`MEM('o011706, 16'o005715);
`MEM('o011710, 16'o001403);
`MEM('o011712, 16'o112720);
`MEM('o011714, 16'o000055);
`MEM('o011716, 16'o000402);
`MEM('o011720, 16'o112720);
`MEM('o011722, 16'o000040);
`MEM('o011724, 16'o062716);
`MEM('o011726, 16'o000060);
`MEM('o011730, 16'o112620);
`MEM('o011732, 16'o005716);
`MEM('o011734, 16'o002373);
`MEM('o011736, 16'o112710);
`MEM('o011740, 16'o000040);
`MEM('o011742, 16'o062706);
`MEM('o011744, 16'o000006);
`MEM('o011746, 16'o012605);
`MEM('o011750, 16'o000207);
`MEM('o011752, 16'o010546);
`MEM('o011754, 16'o010003);
`MEM('o011756, 16'o010105);
`MEM('o011760, 16'o005002);
`MEM('o011762, 16'o005004);
`MEM('o011764, 16'o104462);
`MEM('o011766, 16'o010300);
`MEM('o011770, 16'o010201);
`MEM('o011772, 16'o012605);
`MEM('o011774, 16'o000207);
`MEM('o011776, 16'o005000);
`MEM('o012000, 16'o005001);
`MEM('o012002, 16'o012746);
`MEM('o012004, 16'o000041);
`MEM('o012006, 16'o006000);
`MEM('o012010, 16'o006001);
`MEM('o012012, 16'o006002);
`MEM('o012014, 16'o006003);
`MEM('o012016, 16'o103003);
`MEM('o012020, 16'o060501);
`MEM('o012022, 16'o005500);
`MEM('o012024, 16'o060400);
`MEM('o012026, 16'o005316);
`MEM('o012030, 16'o001366);
`MEM('o012032, 16'o005726);
`MEM('o012034, 16'o000207);
`MEM('o012036, 16'o012746);
`MEM('o012040, 16'o000040);
`MEM('o012042, 16'o010446);
`MEM('o012044, 16'o010546);
`MEM('o012046, 16'o005466);
`MEM('o012050, 16'o000002);
`MEM('o012052, 16'o005416);
`MEM('o012054, 16'o005666);
`MEM('o012056, 16'o000002);
`MEM('o012060, 16'o061601);
`MEM('o012062, 16'o005500);
`MEM('o012064, 16'o066600);
`MEM('o012066, 16'o000002);
`MEM('o012070, 16'o103445);
`MEM('o012072, 16'o005046);
`MEM('o012074, 16'o006103);
`MEM('o012076, 16'o006102);
`MEM('o012100, 16'o006101);
`MEM('o012102, 16'o006100);
`MEM('o012104, 16'o005716);
`MEM('o012106, 16'o001410);
`MEM('o012110, 16'o005016);
`MEM('o012112, 16'o066601);
`MEM('o012114, 16'o000002);
`MEM('o012116, 16'o005500);
`MEM('o012120, 16'o005516);
`MEM('o012122, 16'o066600);
`MEM('o012124, 16'o000004);
`MEM('o012126, 16'o000404);
`MEM('o012130, 16'o060501);
`MEM('o012132, 16'o005500);
`MEM('o012134, 16'o005516);
`MEM('o012136, 16'o060400);
`MEM('o012140, 16'o005516);
`MEM('o012142, 16'o005716);
`MEM('o012144, 16'o001401);
`MEM('o012146, 16'o005203);
`MEM('o012150, 16'o005366);
`MEM('o012152, 16'o000006);
`MEM('o012154, 16'o003347);
`MEM('o012156, 16'o006003);
`MEM('o012160, 16'o103404);
`MEM('o012162, 16'o060501);
`MEM('o012164, 16'o005500);
`MEM('o012166, 16'o060400);
`MEM('o012170, 16'o000241);
`MEM('o012172, 16'o006103);
`MEM('o012174, 16'o062706);
`MEM('o012176, 16'o000010);
`MEM('o012200, 16'o000242);
`MEM('o012202, 16'o000207);
`MEM('o012204, 16'o062706);
`MEM('o012206, 16'o000006);
`MEM('o012210, 16'o104773);
`MEM('o012212, 16'o000262);
`MEM('o012214, 16'o000207);
`MEM('o012216, 16'o010546);
`MEM('o012220, 16'o010046);
`MEM('o012222, 16'o012146);
`MEM('o012224, 16'o012146);
`MEM('o012226, 16'o011146);
`MEM('o012230, 16'o012002);
`MEM('o012232, 16'o012001);
`MEM('o012234, 16'o011000);
`MEM('o012236, 16'o020016);
`MEM('o012240, 16'o101412);
`MEM('o012242, 16'o010604);
`MEM('o012244, 16'o010003);
`MEM('o012246, 16'o011400);
`MEM('o012250, 16'o010324);
`MEM('o012252, 16'o010103);
`MEM('o012254, 16'o011401);
`MEM('o012256, 16'o010324);
`MEM('o012260, 16'o010203);
`MEM('o012262, 16'o011402);
`MEM('o012264, 16'o010324);
`MEM('o012266, 16'o161600);
`MEM('o012270, 16'o001431);
`MEM('o012272, 16'o100003);
`MEM('o012274, 16'o020027);
`MEM('o012276, 16'o177741);
`MEM('o012300, 16'o002005);
`MEM('o012302, 16'o016605);
`MEM('o012304, 16'o000002);
`MEM('o012306, 16'o016603);
`MEM('o012310, 16'o000004);
`MEM('o012312, 16'o000434);
`MEM('o012314, 16'o020027);
`MEM('o012316, 16'o177760);
`MEM('o012320, 16'o003007);
`MEM('o012322, 16'o062700);
`MEM('o012324, 16'o000020);
`MEM('o012326, 16'o010102);
`MEM('o012330, 16'o005001);
`MEM('o012332, 16'o005702);
`MEM('o012334, 16'o100001);
`MEM('o012336, 16'o005101);
`MEM('o012340, 16'o005700);
`MEM('o012342, 16'o001404);
`MEM('o012344, 16'o006201);
`MEM('o012346, 16'o006002);
`MEM('o012350, 16'o005200);
`MEM('o012352, 16'o001374);
`MEM('o012354, 16'o016605);
`MEM('o012356, 16'o000002);
`MEM('o012360, 16'o016603);
`MEM('o012362, 16'o000004);
`MEM('o012364, 16'o060203);
`MEM('o012366, 16'o005505);
`MEM('o012370, 16'o102421);
`MEM('o012372, 16'o060105);
`MEM('o012374, 16'o102003);
`MEM('o012376, 16'o006005);
`MEM('o012400, 16'o006003);
`MEM('o012402, 16'o005216);
`MEM('o012404, 16'o016600);
`MEM('o012406, 16'o000006);
`MEM('o012410, 16'o010001);
`MEM('o012412, 16'o010320);
`MEM('o012414, 16'o010520);
`MEM('o012416, 16'o011620);
`MEM('o012420, 16'o010100);
`MEM('o012422, 16'o062706);
`MEM('o012424, 16'o000010);
`MEM('o012426, 16'o012605);
`MEM('o012430, 16'o000167);
`MEM('o012432, 16'o000546);
`MEM('o012434, 16'o060105);
`MEM('o012436, 16'o103762);
`MEM('o012440, 16'o000756);
`MEM('o012442, 16'o010004);
`MEM('o012444, 16'o162706);
`MEM('o012446, 16'o000006);
`MEM('o012450, 16'o010600);
`MEM('o012452, 16'o104424);
`MEM('o012454, 16'o010400);
`MEM('o012456, 16'o010601);
`MEM('o012460, 16'o104420);
`MEM('o012462, 16'o062706);
`MEM('o012464, 16'o000006);
`MEM('o012466, 16'o000207);
`MEM('o012470, 16'o104432);
`MEM('o012472, 16'o005761);
`MEM('o012474, 16'o000002);
`MEM('o012476, 16'o002010);
`MEM('o012500, 16'o012102);
`MEM('o012502, 16'o012103);
`MEM('o012504, 16'o005403);
`MEM('o012506, 16'o005402);
`MEM('o012510, 16'o005603);
`MEM('o012512, 16'o010220);
`MEM('o012514, 16'o010320);
`MEM('o012516, 16'o012120);
`MEM('o012520, 16'o000207);
`MEM('o012522, 16'o104432);
`MEM('o012524, 16'o012701);
`MEM('o012526, 16'o010666);
`MEM('o012530, 16'o005760);
`MEM('o012532, 16'o000002);
`MEM('o012534, 16'o003003);
`MEM('o012536, 16'o001403);
`MEM('o012540, 16'o104424);
`MEM('o012542, 16'o000207);
`MEM('o012544, 16'o104432);
`MEM('o012546, 16'o000207);
`MEM('o012550, 16'o010546);
`MEM('o012552, 16'o010046);
`MEM('o012554, 16'o005046);
`MEM('o012556, 16'o012105);
`MEM('o012560, 16'o012104);
`MEM('o012562, 16'o005704);
`MEM('o012564, 16'o001477);
`MEM('o012566, 16'o002004);
`MEM('o012570, 16'o005404);
`MEM('o012572, 16'o005405);
`MEM('o012574, 16'o005604);
`MEM('o012576, 16'o005216);
`MEM('o012600, 16'o012003);
`MEM('o012602, 16'o012002);
`MEM('o012604, 16'o001563);
`MEM('o012606, 16'o003004);
`MEM('o012610, 16'o005402);
`MEM('o012612, 16'o005403);
`MEM('o012614, 16'o005602);
`MEM('o012616, 16'o005316);
`MEM('o012620, 16'o011101);
`MEM('o012622, 16'o005401);
`MEM('o012624, 16'o061001);
`MEM('o012626, 16'o006001);
`MEM('o012630, 16'o006101);
`MEM('o012632, 16'o102054);
`MEM('o012634, 16'o062701);
`MEM('o012636, 16'o100000);
`MEM('o012640, 16'o010146);
`MEM('o012642, 16'o010301);
`MEM('o012644, 16'o010200);
`MEM('o012646, 16'o005002);
`MEM('o012650, 16'o005003);
`MEM('o012652, 16'o006000);
`MEM('o012654, 16'o006001);
`MEM('o012656, 16'o006002);
`MEM('o012660, 16'o104464);
`MEM('o012662, 16'o005404);
`MEM('o012664, 16'o005405);
`MEM('o012666, 16'o005604);
`MEM('o012670, 16'o006301);
`MEM('o012672, 16'o006100);
`MEM('o012674, 16'o060501);
`MEM('o012676, 16'o005500);
`MEM('o012700, 16'o060400);
`MEM('o012702, 16'o002403);
`MEM('o012704, 16'o062703);
`MEM('o012706, 16'o000001);
`MEM('o012710, 16'o005502);
`MEM('o012712, 16'o000241);
`MEM('o012714, 16'o006002);
`MEM('o012716, 16'o006003);
`MEM('o012720, 16'o005216);
`MEM('o012722, 16'o005766);
`MEM('o012724, 16'o000002);
`MEM('o012726, 16'o001403);
`MEM('o012730, 16'o005402);
`MEM('o012732, 16'o005403);
`MEM('o012734, 16'o005602);
`MEM('o012736, 16'o016600);
`MEM('o012740, 16'o000004);
`MEM('o012742, 16'o010320);
`MEM('o012744, 16'o010220);
`MEM('o012746, 16'o012610);
`MEM('o012750, 16'o022626);
`MEM('o012752, 16'o012605);
`MEM('o012754, 16'o024040);
`MEM('o012756, 16'o010001);
`MEM('o012760, 16'o000167);
`MEM('o012762, 16'o000216);
`MEM('o012764, 16'o022626);
`MEM('o012766, 16'o104773);
`MEM('o012770, 16'o012605);
`MEM('o012772, 16'o000262);
`MEM('o012774, 16'o000207);
`MEM('o012776, 16'o010546);
`MEM('o013000, 16'o010046);
`MEM('o013002, 16'o012105);
`MEM('o013004, 16'o012104);
`MEM('o013006, 16'o011101);
`MEM('o013010, 16'o005046);
`MEM('o013012, 16'o005704);
`MEM('o013014, 16'o001457);
`MEM('o013016, 16'o100004);
`MEM('o013020, 16'o005404);
`MEM('o013022, 16'o005405);
`MEM('o013024, 16'o005604);
`MEM('o013026, 16'o005316);
`MEM('o013030, 16'o012003);
`MEM('o013032, 16'o012002);
`MEM('o013034, 16'o001447);
`MEM('o013036, 16'o100004);
`MEM('o013040, 16'o005402);
`MEM('o013042, 16'o005403);
`MEM('o013044, 16'o005602);
`MEM('o013046, 16'o005216);
`MEM('o013050, 16'o061001);
`MEM('o013052, 16'o006001);
`MEM('o013054, 16'o006101);
`MEM('o013056, 16'o102342);
`MEM('o013060, 16'o062701);
`MEM('o013062, 16'o100000);
`MEM('o013064, 16'o010146);
`MEM('o013066, 16'o104462);
`MEM('o013070, 16'o005216);
`MEM('o013072, 16'o006102);
`MEM('o013074, 16'o006101);
`MEM('o013076, 16'o006100);
`MEM('o013100, 16'o102402);
`MEM('o013102, 16'o005316);
`MEM('o013104, 16'o000772);
`MEM('o013106, 16'o006000);
`MEM('o013110, 16'o006001);
`MEM('o013112, 16'o005501);
`MEM('o013114, 16'o005500);
`MEM('o013116, 16'o102002);
`MEM('o013120, 16'o005216);
`MEM('o013122, 16'o000771);
`MEM('o013124, 16'o012602);
`MEM('o013126, 16'o005726);
`MEM('o013130, 16'o001403);
`MEM('o013132, 16'o005400);
`MEM('o013134, 16'o005401);
`MEM('o013136, 16'o005600);
`MEM('o013140, 16'o012603);
`MEM('o013142, 16'o010123);
`MEM('o013144, 16'o010023);
`MEM('o013146, 16'o010213);
`MEM('o013150, 16'o012605);
`MEM('o013152, 16'o000207);
`MEM('o013154, 16'o005000);
`MEM('o013156, 16'o005001);
`MEM('o013160, 16'o005002);
`MEM('o013162, 16'o005726);
`MEM('o013164, 16'o000765);
`MEM('o013166, 16'o005020);
`MEM('o013170, 16'o010120);
`MEM('o013172, 16'o012710);
`MEM('o013174, 16'o100017);
`MEM('o013176, 16'o024040);
`MEM('o013200, 16'o010001);
`MEM('o013202, 16'o012104);
`MEM('o013204, 16'o012102);
`MEM('o013206, 16'o012103);
`MEM('o013210, 16'o010301);
`MEM('o013212, 16'o005702);
`MEM('o013214, 16'o001004);
`MEM('o013216, 16'o005704);
`MEM('o013220, 16'o001002);
`MEM('o013222, 16'o005003);
`MEM('o013224, 16'o000420);
`MEM('o013226, 16'o005203);
`MEM('o013230, 16'o005303);
`MEM('o013232, 16'o006304);
`MEM('o013234, 16'o006102);
`MEM('o013236, 16'o102374);
`MEM('o013240, 16'o103010);
`MEM('o013242, 16'o001007);
`MEM('o013244, 16'o005704);
`MEM('o013246, 16'o001004);
`MEM('o013250, 16'o000261);
`MEM('o013252, 16'o006002);
`MEM('o013254, 16'o005203);
`MEM('o013256, 16'o005201);
`MEM('o013260, 16'o000261);
`MEM('o013262, 16'o006002);
`MEM('o013264, 16'o006004);
`MEM('o013266, 16'o010420);
`MEM('o013270, 16'o010220);
`MEM('o013272, 16'o010320);
`MEM('o013274, 16'o020301);
`MEM('o013276, 16'o101002);
`MEM('o013300, 16'o000242);
`MEM('o013302, 16'o000207);
`MEM('o013304, 16'o000262);
`MEM('o013306, 16'o000207);
`MEM('o013310, 16'o010102);
`MEM('o013312, 16'o010004);
`MEM('o013314, 16'o012224);
`MEM('o013316, 16'o012224);
`MEM('o013320, 16'o012224);
`MEM('o013322, 16'o000207);
`MEM('o013324, 16'o010146);
`MEM('o013326, 16'o104454);
`MEM('o013330, 16'o010600);
`MEM('o013332, 16'o016601);
`MEM('o013334, 16'o000006);
`MEM('o013336, 16'o104422);
`MEM('o013340, 16'o016601);
`MEM('o013342, 16'o000002);
`MEM('o013344, 16'o062706);
`MEM('o013346, 16'o000010);
`MEM('o013350, 16'o005401);
`MEM('o013352, 16'o000207);
`MEM('o013354, 16'o012602);
`MEM('o013356, 16'o062700);
`MEM('o013360, 16'o000006);
`MEM('o013362, 16'o014046);
`MEM('o013364, 16'o014046);
`MEM('o013366, 16'o014046);
`MEM('o013370, 16'o010207);
`MEM('o013372, 16'o012103);
`MEM('o013374, 16'o012102);
`MEM('o013376, 16'o011104);
`MEM('o013400, 16'o100021);
`MEM('o013402, 16'o024141);
`MEM('o013404, 16'o020427);
`MEM('o013406, 16'o100037);
`MEM('o013410, 16'o103337);
`MEM('o013412, 16'o162704);
`MEM('o013414, 16'o100037);
`MEM('o013416, 16'o006202);
`MEM('o013420, 16'o006003);
`MEM('o013422, 16'o005204);
`MEM('o013424, 16'o002774);
`MEM('o013426, 16'o010001);
`MEM('o013430, 16'o010320);
`MEM('o013432, 16'o010220);
`MEM('o013434, 16'o012710);
`MEM('o013436, 16'o100037);
`MEM('o013440, 16'o010100);
`MEM('o013442, 16'o000657);
`MEM('o013444, 16'o005702);
`MEM('o013446, 16'o100004);
`MEM('o013450, 16'o012701);
`MEM('o013452, 16'o010666);
`MEM('o013454, 16'o000167);
`MEM('o013456, 16'o177020);
`MEM('o013460, 16'o005020);
`MEM('o013462, 16'o005020);
`MEM('o013464, 16'o005010);
`MEM('o013466, 16'o000207);
`MEM('o013470, 16'o012102);
`MEM('o013472, 16'o012103);
`MEM('o013474, 16'o011104);
`MEM('o013476, 16'o020427);
`MEM('o013500, 16'o100017);
`MEM('o013502, 16'o101013);
`MEM('o013504, 16'o001410);
`MEM('o013506, 16'o020427);
`MEM('o013510, 16'o100000);
`MEM('o013512, 16'o103410);
`MEM('o013514, 16'o162704);
`MEM('o013516, 16'o100017);
`MEM('o013520, 16'o006203);
`MEM('o013522, 16'o005204);
`MEM('o013524, 16'o001375);
`MEM('o013526, 16'o010300);
`MEM('o013530, 16'o000207);
`MEM('o013532, 16'o104771);
`MEM('o013534, 16'o005000);
`MEM('o013536, 16'o000207);
`MEM('o013540, 16'o042120);
`MEM('o013542, 16'o026520);
`MEM('o013544, 16'o030461);
`MEM('o013546, 16'o041040);
`MEM('o013550, 16'o051501);
`MEM('o013552, 16'o041511);
`MEM('o013554, 16'o020054);
`MEM('o013556, 16'o042526);
`MEM('o013560, 16'o051522);
`MEM('o013562, 16'o047511);
`MEM('o013564, 16'o020116);
`MEM('o013566, 16'o030060);
`MEM('o013570, 16'o040467);
`MEM('o013572, 16'o005015);
`MEM('o013574, 16'o047452);
`MEM('o013576, 16'o000040);
`MEM('o013600, 16'o000000);
`MEM('o013602, 16'o000000);
`MEM('o013604, 16'o000000);
`MEM('o013606, 16'o000000);
`MEM('o013610, 16'o000000);
`MEM('o013612, 16'o000000);
`MEM('o013614, 16'o000000);
`MEM('o013616, 16'o000000);
`MEM('o013620, 16'o000000);
`MEM('o013622, 16'o000000);
`MEM('o013624, 16'o000000);
`MEM('o013626, 16'o000000);
`MEM('o013630, 16'o000000);
`MEM('o013632, 16'o000000);
`MEM('o013634, 16'o000000);
`MEM('o013636, 16'o000000);
`MEM('o013640, 16'o000000);
`MEM('o013642, 16'o000000);
`MEM('o013644, 16'o000000);
`MEM('o013646, 16'o000000);
`MEM('o013650, 16'o077474);
`MEM('o013652, 16'o000354);
`MEM('o013654, 16'o017016);
`MEM('o013656, 16'o016170);
`MEM('o013660, 16'o000000);
`MEM('o013662, 16'o000000);
`MEM('o013664, 16'o000000);
`MEM('o013666, 16'o000000);
`MEM('o013670, 16'o000000);
`MEM('o013672, 16'o000037);
`MEM('o013674, 16'o000000);
`MEM('o013676, 16'o000000);
`MEM('o013700, 16'o000001);
`MEM('o013702, 16'o000000);
`MEM('o013704, 16'o000000);
`MEM('o013706, 16'o000000);
`MEM('o013710, 16'o030355);
`MEM('o013712, 16'o013660);
`MEM('o013714, 16'o010146);
`MEM('o013716, 16'o010046);
`MEM('o013720, 16'o162706);
`MEM('o013722, 16'o000006);
`MEM('o013724, 16'o010001);
`MEM('o013726, 16'o010600);
`MEM('o013730, 16'o004767);
`MEM('o013732, 16'o000030);
`MEM('o013734, 16'o016601);
`MEM('o013736, 16'o000010);
`MEM('o013740, 16'o010600);
`MEM('o013742, 16'o104430);
`MEM('o013744, 16'o016600);
`MEM('o013746, 16'o000006);
`MEM('o013750, 16'o010601);
`MEM('o013752, 16'o004767);
`MEM('o013754, 16'o000302);
`MEM('o013756, 16'o062706);
`MEM('o013760, 16'o000012);
`MEM('o013762, 16'o000207);
`MEM('o013764, 16'o104456);
`MEM('o013766, 16'o005760);
`MEM('o013770, 16'o000002);
`MEM('o013772, 16'o003004);
`MEM('o013774, 16'o104777);
`MEM('o013776, 16'o062706);
`MEM('o014000, 16'o000004);
`MEM('o014002, 16'o000207);
`MEM('o014004, 16'o010001);
`MEM('o014006, 16'o005721);
`MEM('o014010, 16'o001014);
`MEM('o014012, 16'o022127);
`MEM('o014014, 16'o040000);
`MEM('o014016, 16'o001011);
`MEM('o014020, 16'o022127);
`MEM('o014022, 16'o100001);
`MEM('o014024, 16'o001006);
`MEM('o014026, 16'o005020);
`MEM('o014030, 16'o005020);
`MEM('o014032, 16'o005020);
`MEM('o014034, 16'o062706);
`MEM('o014036, 16'o000004);
`MEM('o014040, 16'o000207);
`MEM('o014042, 16'o016046);
`MEM('o014044, 16'o000004);
`MEM('o014046, 16'o062716);
`MEM('o014050, 16'o100000);
`MEM('o014052, 16'o012760);
`MEM('o014054, 16'o100000);
`MEM('o014056, 16'o000004);
`MEM('o014060, 16'o011601);
`MEM('o014062, 16'o162706);
`MEM('o014064, 16'o000006);
`MEM('o014066, 16'o010600);
`MEM('o014070, 16'o104436);
`MEM('o014072, 16'o016600);
`MEM('o014074, 16'o000010);
`MEM('o014076, 16'o104454);
`MEM('o014100, 16'o012701);
`MEM('o014102, 16'o014214);
`MEM('o014104, 16'o104422);
`MEM('o014106, 16'o010600);
`MEM('o014110, 16'o012701);
`MEM('o014112, 16'o014214);
`MEM('o014114, 16'o104420);
`MEM('o014116, 16'o016600);
`MEM('o014120, 16'o000016);
`MEM('o014122, 16'o010601);
`MEM('o014124, 16'o104426);
`MEM('o014126, 16'o012704);
`MEM('o014130, 16'o014230);
`MEM('o014132, 16'o016600);
`MEM('o014134, 16'o000016);
`MEM('o014136, 16'o012703);
`MEM('o014140, 16'o000004);
`MEM('o014142, 16'o104450);
`MEM('o014144, 16'o104452);
`MEM('o014146, 16'o016600);
`MEM('o014150, 16'o000016);
`MEM('o014152, 16'o012701);
`MEM('o014154, 16'o014506);
`MEM('o014156, 16'o104422);
`MEM('o014160, 16'o062706);
`MEM('o014162, 16'o000006);
`MEM('o014164, 16'o010600);
`MEM('o014166, 16'o012701);
`MEM('o014170, 16'o014222);
`MEM('o014172, 16'o104430);
`MEM('o014174, 16'o010601);
`MEM('o014176, 16'o016600);
`MEM('o014200, 16'o000010);
`MEM('o014202, 16'o104420);
`MEM('o014204, 16'o062706);
`MEM('o014206, 16'o000014);
`MEM('o014210, 16'o000242);
`MEM('o014212, 16'o000207);
`MEM('o014214, 16'o074626);
`MEM('o014216, 16'o055202);
`MEM('o014220, 16'o100000);
`MEM('o014222, 16'o005776);
`MEM('o014224, 16'o054271);
`MEM('o014226, 16'o100000);
`MEM('o014230, 16'o125112);
`MEM('o014232, 16'o046414);
`MEM('o014234, 16'o077777);
`MEM('o014236, 16'o007411);
`MEM('o014240, 16'o063120);
`MEM('o014242, 16'o077777);
`MEM('o014244, 16'o066333);
`MEM('o014246, 16'o052525);
`MEM('o014250, 16'o100000);
`MEM('o014252, 16'o177772);
`MEM('o014254, 16'o077777);
`MEM('o014256, 16'o100001);
`MEM('o014260, 16'o104456);
`MEM('o014262, 16'o026027);
`MEM('o014264, 16'o000004);
`MEM('o014266, 16'o100016);
`MEM('o014270, 16'o101241);
`MEM('o014272, 16'o012701);
`MEM('o014274, 16'o014500);
`MEM('o014276, 16'o104446);
`MEM('o014300, 16'o016600);
`MEM('o014302, 16'o000002);
`MEM('o014304, 16'o012701);
`MEM('o014306, 16'o014506);
`MEM('o014310, 16'o104430);
`MEM('o014312, 16'o016600);
`MEM('o014314, 16'o000002);
`MEM('o014316, 16'o104454);
`MEM('o014320, 16'o104454);
`MEM('o014322, 16'o010600);
`MEM('o014324, 16'o012701);
`MEM('o014326, 16'o014514);
`MEM('o014330, 16'o104420);
`MEM('o014332, 16'o010600);
`MEM('o014334, 16'o010001);
`MEM('o014336, 16'o104424);
`MEM('o014340, 16'o005266);
`MEM('o014342, 16'o000012);
`MEM('o014344, 16'o016600);
`MEM('o014346, 16'o000016);
`MEM('o014350, 16'o010001);
`MEM('o014352, 16'o104430);
`MEM('o014354, 16'o016600);
`MEM('o014356, 16'o000016);
`MEM('o014360, 16'o012701);
`MEM('o014362, 16'o014530);
`MEM('o014364, 16'o104420);
`MEM('o014366, 16'o012700);
`MEM('o014370, 16'o014522);
`MEM('o014372, 16'o104454);
`MEM('o014374, 16'o010600);
`MEM('o014376, 16'o016601);
`MEM('o014400, 16'o000024);
`MEM('o014402, 16'o104426);
`MEM('o014404, 16'o010600);
`MEM('o014406, 16'o010001);
`MEM('o014410, 16'o062701);
`MEM('o014412, 16'o000006);
`MEM('o014414, 16'o104420);
`MEM('o014416, 16'o010601);
`MEM('o014420, 16'o010100);
`MEM('o014422, 16'o062700);
`MEM('o014424, 16'o000014);
`MEM('o014426, 16'o104426);
`MEM('o014430, 16'o062706);
`MEM('o014432, 16'o000014);
`MEM('o014434, 16'o010600);
`MEM('o014436, 16'o012701);
`MEM('o014440, 16'o010666);
`MEM('o014442, 16'o104420);
`MEM('o014444, 16'o010600);
`MEM('o014446, 16'o010001);
`MEM('o014450, 16'o104430);
`MEM('o014452, 16'o010601);
`MEM('o014454, 16'o016600);
`MEM('o014456, 16'o000010);
`MEM('o014460, 16'o104432);
`MEM('o014462, 16'o016600);
`MEM('o014464, 16'o000010);
`MEM('o014466, 16'o066660);
`MEM('o014470, 16'o000006);
`MEM('o014472, 16'o000004);
`MEM('o014474, 16'o000167);
`MEM('o014476, 16'o177504);
`MEM('o014500, 16'o016624);
`MEM('o014502, 16'o056125);
`MEM('o014504, 16'o100001);
`MEM('o014506, 16'o005776);
`MEM('o014510, 16'o054271);
`MEM('o014512, 16'o077777);
`MEM('o014514, 16'o037347);
`MEM('o014516, 16'o117741);
`MEM('o014520, 16'o100004);
`MEM('o014522, 16'o041565);
`MEM('o014524, 16'o132306);
`MEM('o014526, 16'o100012);
`MEM('o014530, 16'o026570);
`MEM('o014532, 16'o074056);
`MEM('o014534, 16'o100006);
`MEM('o014536, 16'o162766);
`MEM('o014540, 16'o000002);
`MEM('o014542, 16'o000002);
`MEM('o014544, 16'o016600);
`MEM('o014546, 16'o000010);
`MEM('o014550, 16'o016601);
`MEM('o014552, 16'o000012);
`MEM('o014554, 16'o010046);
`MEM('o014556, 16'o104430);
`MEM('o014560, 16'o062766);
`MEM('o014562, 16'o000006);
`MEM('o014564, 16'o000014);
`MEM('o014566, 16'o011600);
`MEM('o014570, 16'o016601);
`MEM('o014572, 16'o000014);
`MEM('o014574, 16'o104420);
`MEM('o014576, 16'o005766);
`MEM('o014600, 16'o000004);
`MEM('o014602, 16'o001407);
`MEM('o014604, 16'o011600);
`MEM('o014606, 16'o016601);
`MEM('o014610, 16'o000010);
`MEM('o014612, 16'o104430);
`MEM('o014614, 16'o005366);
`MEM('o014616, 16'o000004);
`MEM('o014620, 16'o000757);
`MEM('o014622, 16'o011600);
`MEM('o014624, 16'o016601);
`MEM('o014626, 16'o000006);
`MEM('o014630, 16'o104430);
`MEM('o014632, 16'o005726);
`MEM('o014634, 16'o012603);
`MEM('o014636, 16'o062706);
`MEM('o014640, 16'o000026);
`MEM('o014642, 16'o010346);
`MEM('o014644, 16'o000207);
`MEM('o014646, 16'o012603);
`MEM('o014650, 16'o005046);
`MEM('o014652, 16'o010146);
`MEM('o014654, 16'o010046);
`MEM('o014656, 16'o104432);
`MEM('o014660, 16'o010307);
`MEM('o014662, 16'o012603);
`MEM('o014664, 16'o000772);
`MEM('o014666, 16'o012601);
`MEM('o014670, 16'o104454);
`MEM('o014672, 16'o010146);
`MEM('o014674, 16'o010446);
`MEM('o014676, 16'o010346);
`MEM('o014700, 16'o010046);
`MEM('o014702, 16'o010001);
`MEM('o014704, 16'o104430);
`MEM('o014706, 16'o012600);
`MEM('o014710, 16'o012603);
`MEM('o014712, 16'o012604);
`MEM('o014714, 16'o012601);
`MEM('o014716, 16'o104454);
`MEM('o014720, 16'o010446);
`MEM('o014722, 16'o010046);
`MEM('o014724, 16'o010646);
`MEM('o014726, 16'o062716);
`MEM('o014730, 16'o000006);
`MEM('o014732, 16'o010646);
`MEM('o014734, 16'o062716);
`MEM('o014736, 16'o000016);
`MEM('o014740, 16'o010346);
`MEM('o014742, 16'o010107);
`MEM('o014744, 16'o016600);
`MEM('o014746, 16'o000002);
`MEM('o014750, 16'o104430);
`MEM('o014752, 16'o012666);
`MEM('o014754, 16'o000002);
`MEM('o014756, 16'o011601);
`MEM('o014760, 16'o104442);
`MEM('o014762, 16'o010046);
`MEM('o014764, 16'o011601);
`MEM('o014766, 16'o162706);
`MEM('o014770, 16'o000006);
`MEM('o014772, 16'o010600);
`MEM('o014774, 16'o104436);
`MEM('o014776, 16'o010601);
`MEM('o015000, 16'o016600);
`MEM('o015002, 16'o000010);
`MEM('o015004, 16'o104422);
`MEM('o015006, 16'o062706);
`MEM('o015010, 16'o000006);
`MEM('o015012, 16'o016646);
`MEM('o015014, 16'o000004);
`MEM('o015016, 16'o000207);
`MEM('o015020, 16'o104444);
`MEM('o015022, 16'o005760);
`MEM('o015024, 16'o000002);
`MEM('o015026, 16'o002005);
`MEM('o015030, 16'o010001);
`MEM('o015032, 16'o104424);
`MEM('o015034, 16'o005266);
`MEM('o015036, 16'o000004);
`MEM('o015040, 16'o000404);
`MEM('o015042, 16'o001003);
`MEM('o015044, 16'o062706);
`MEM('o015046, 16'o000006);
`MEM('o015050, 16'o000207);
`MEM('o015052, 16'o012701);
`MEM('o015054, 16'o015206);
`MEM('o015056, 16'o104446);
`MEM('o015060, 16'o012602);
`MEM('o015062, 16'o042702);
`MEM('o015064, 16'o177774);
`MEM('o015066, 16'o006302);
`MEM('o015070, 16'o062702);
`MEM('o015072, 16'o015176);
`MEM('o015074, 16'o011207);
`MEM('o015076, 16'o012701);
`MEM('o015100, 16'o010666);
`MEM('o015102, 16'o011600);
`MEM('o015104, 16'o104422);
`MEM('o015106, 16'o011600);
`MEM('o015110, 16'o010001);
`MEM('o015112, 16'o104424);
`MEM('o015114, 16'o000404);
`MEM('o015116, 16'o012701);
`MEM('o015120, 16'o010666);
`MEM('o015122, 16'o011600);
`MEM('o015124, 16'o104422);
`MEM('o015126, 16'o011600);
`MEM('o015130, 16'o012704);
`MEM('o015132, 16'o015214);
`MEM('o015134, 16'o012703);
`MEM('o015136, 16'o000006);
`MEM('o015140, 16'o104450);
`MEM('o015142, 16'o104452);
`MEM('o015144, 16'o005766);
`MEM('o015146, 16'o000004);
`MEM('o015150, 16'o001735);
`MEM('o015152, 16'o011600);
`MEM('o015154, 16'o010001);
`MEM('o015156, 16'o104424);
`MEM('o015160, 16'o000731);
`MEM('o015162, 16'o104444);
`MEM('o015164, 16'o012701);
`MEM('o015166, 16'o015252);
`MEM('o015170, 16'o104420);
`MEM('o015172, 16'o011600);
`MEM('o015174, 16'o000712);
`MEM('o015176, 16'o015126);
`MEM('o015200, 16'o015076);
`MEM('o015202, 16'o015106);
`MEM('o015204, 16'o015116);
`MEM('o015206, 16'o140671);
`MEM('o015210, 16'o050574);
`MEM('o015212, 16'o100000);
`MEM('o015214, 16'o017676);
`MEM('o015216, 16'o106516);
`MEM('o015220, 16'o077756);
`MEM('o015222, 16'o175316);
`MEM('o015224, 16'o051777);
`MEM('o015226, 16'o077764);
`MEM('o015230, 16'o156214);
`MEM('o015232, 16'o131513);
`MEM('o015234, 16'o077771);
`MEM('o015236, 16'o167376);
`MEM('o015240, 16'o050632);
`MEM('o015242, 16'o077775);
`MEM('o015244, 16'o006165);
`MEM('o015246, 16'o126521);
`MEM('o015250, 16'o100000);
`MEM('o015252, 16'o166516);
`MEM('o015254, 16'o062207);
`MEM('o015256, 16'o100001);
`MEM('o015260, 16'o005046);
`MEM('o015262, 16'o104444);
`MEM('o015264, 16'o005760);
`MEM('o015266, 16'o000002);
`MEM('o015270, 16'o001530);
`MEM('o015272, 16'o002004);
`MEM('o015274, 16'o005266);
`MEM('o015276, 16'o000006);
`MEM('o015300, 16'o010001);
`MEM('o015302, 16'o104424);
`MEM('o015304, 16'o012701);
`MEM('o015306, 16'o010666);
`MEM('o015310, 16'o011600);
`MEM('o015312, 16'o104434);
`MEM('o015314, 16'o002017);
`MEM('o015316, 16'o005266);
`MEM('o015320, 16'o000004);
`MEM('o015322, 16'o012700);
`MEM('o015324, 16'o010666);
`MEM('o015326, 16'o104454);
`MEM('o015330, 16'o010600);
`MEM('o015332, 16'o016601);
`MEM('o015334, 16'o000006);
`MEM('o015336, 16'o104426);
`MEM('o015340, 16'o010601);
`MEM('o015342, 16'o016600);
`MEM('o015344, 16'o000006);
`MEM('o015346, 16'o104432);
`MEM('o015350, 16'o062706);
`MEM('o015352, 16'o000006);
`MEM('o015354, 16'o012701);
`MEM('o015356, 16'o015562);
`MEM('o015360, 16'o011600);
`MEM('o015362, 16'o104434);
`MEM('o015364, 16'o003404);
`MEM('o015366, 16'o005046);
`MEM('o015370, 16'o005046);
`MEM('o015372, 16'o005046);
`MEM('o015374, 16'o000430);
`MEM('o015376, 16'o012700);
`MEM('o015400, 16'o015576);
`MEM('o015402, 16'o104454);
`MEM('o015404, 16'o016600);
`MEM('o015406, 16'o000006);
`MEM('o015410, 16'o104454);
`MEM('o015412, 16'o012701);
`MEM('o015414, 16'o015570);
`MEM('o015416, 16'o104430);
`MEM('o015420, 16'o016600);
`MEM('o015422, 16'o000014);
`MEM('o015424, 16'o012701);
`MEM('o015426, 16'o010666);
`MEM('o015430, 16'o104422);
`MEM('o015432, 16'o010600);
`MEM('o015434, 16'o012701);
`MEM('o015436, 16'o015570);
`MEM('o015440, 16'o104420);
`MEM('o015442, 16'o016600);
`MEM('o015444, 16'o000014);
`MEM('o015446, 16'o010601);
`MEM('o015450, 16'o104426);
`MEM('o015452, 16'o062706);
`MEM('o015454, 16'o000006);
`MEM('o015456, 16'o016600);
`MEM('o015460, 16'o000006);
`MEM('o015462, 16'o012704);
`MEM('o015464, 16'o015604);
`MEM('o015466, 16'o012703);
`MEM('o015470, 16'o000005);
`MEM('o015472, 16'o104450);
`MEM('o015474, 16'o104452);
`MEM('o015476, 16'o010601);
`MEM('o015500, 16'o016600);
`MEM('o015502, 16'o000006);
`MEM('o015504, 16'o104420);
`MEM('o015506, 16'o062706);
`MEM('o015510, 16'o000006);
`MEM('o015512, 16'o005766);
`MEM('o015514, 16'o000004);
`MEM('o015516, 16'o001407);
`MEM('o015520, 16'o011600);
`MEM('o015522, 16'o012701);
`MEM('o015524, 16'o015252);
`MEM('o015526, 16'o104422);
`MEM('o015530, 16'o011600);
`MEM('o015532, 16'o010001);
`MEM('o015534, 16'o104424);
`MEM('o015536, 16'o005766);
`MEM('o015540, 16'o000006);
`MEM('o015542, 16'o001403);
`MEM('o015544, 16'o011600);
`MEM('o015546, 16'o010001);
`MEM('o015550, 16'o104424);
`MEM('o015552, 16'o062706);
`MEM('o015554, 16'o000010);
`MEM('o015556, 16'o000242);
`MEM('o015560, 16'o000207);
`MEM('o015562, 16'o050574);
`MEM('o015564, 16'o042230);
`MEM('o015566, 16'o077777);
`MEM('o015570, 16'o165640);
`MEM('o015572, 16'o067331);
`MEM('o015574, 16'o100001);
`MEM('o015576, 16'o044336);
`MEM('o015600, 16'o041405);
`MEM('o015602, 16'o100000);
`MEM('o015604, 16'o113440);
`MEM('o015606, 16'o060462);
`MEM('o015610, 16'o077775);
`MEM('o015612, 16'o107717);
`MEM('o015614, 16'o133556);
`MEM('o015616, 16'o077776);
`MEM('o015620, 16'o155646);
`MEM('o015622, 16'o063141);
`MEM('o015624, 16'o077776);
`MEM('o015626, 16'o131012);
`MEM('o015630, 16'o125252);
`MEM('o015632, 16'o077777);
`MEM('o015634, 16'o177776);
`MEM('o015636, 16'o077777);
`MEM('o015640, 16'o100000);
`MEM('o015642, 16'o104444);
`MEM('o015644, 16'o005760);
`MEM('o015646, 16'o000002);
`MEM('o015650, 16'o001456);
`MEM('o015652, 16'o002004);
`MEM('o015654, 16'o005266);
`MEM('o015656, 16'o000004);
`MEM('o015660, 16'o010001);
`MEM('o015662, 16'o104424);
`MEM('o015664, 16'o005066);
`MEM('o015666, 16'o000002);
`MEM('o015670, 16'o011600);
`MEM('o015672, 16'o022020);
`MEM('o015674, 16'o062710);
`MEM('o015676, 16'o100000);
`MEM('o015700, 16'o006210);
`MEM('o015702, 16'o005566);
`MEM('o015704, 16'o000002);
`MEM('o015706, 16'o011046);
`MEM('o015710, 16'o012710);
`MEM('o015712, 16'o100000);
`MEM('o015714, 16'o016600);
`MEM('o015716, 16'o000002);
`MEM('o015720, 16'o104454);
`MEM('o015722, 16'o012701);
`MEM('o015724, 16'o016076);
`MEM('o015726, 16'o104430);
`MEM('o015730, 16'o016600);
`MEM('o015732, 16'o000010);
`MEM('o015734, 16'o012701);
`MEM('o015736, 16'o016070);
`MEM('o015740, 16'o104420);
`MEM('o015742, 16'o104460);
`MEM('o015744, 16'o104460);
`MEM('o015746, 16'o104460);
`MEM('o015750, 16'o066660);
`MEM('o015752, 16'o000006);
`MEM('o015754, 16'o000004);
`MEM('o015756, 16'o062706);
`MEM('o015760, 16'o000010);
`MEM('o015762, 16'o005766);
`MEM('o015764, 16'o000002);
`MEM('o015766, 16'o001403);
`MEM('o015770, 16'o012701);
`MEM('o015772, 16'o016062);
`MEM('o015774, 16'o104430);
`MEM('o015776, 16'o005766);
`MEM('o016000, 16'o000004);
`MEM('o016002, 16'o001401);
`MEM('o016004, 16'o104775);
`MEM('o016006, 16'o062706);
`MEM('o016010, 16'o000006);
`MEM('o016012, 16'o000242);
`MEM('o016014, 16'o000207);
`MEM('o016016, 16'o010600);
`MEM('o016020, 16'o005720);
`MEM('o016022, 16'o104454);
`MEM('o016024, 16'o010600);
`MEM('o016026, 16'o016601);
`MEM('o016030, 16'o000020);
`MEM('o016032, 16'o104426);
`MEM('o016034, 16'o010601);
`MEM('o016036, 16'o016600);
`MEM('o016040, 16'o000020);
`MEM('o016042, 16'o104420);
`MEM('o016044, 16'o016600);
`MEM('o016046, 16'o000020);
`MEM('o016050, 16'o005360);
`MEM('o016052, 16'o000004);
`MEM('o016054, 16'o062706);
`MEM('o016056, 16'o000006);
`MEM('o016060, 16'o000207);
`MEM('o016062, 16'o074626);
`MEM('o016064, 16'o055202);
`MEM('o016066, 16'o100001);
`MEM('o016070, 16'o125672);
`MEM('o016072, 16'o065324);
`MEM('o016074, 16'o077777);
`MEM('o016076, 16'o067102);
`MEM('o016100, 16'o045612);
`MEM('o016102, 16'o100000);
`MEM('o016104, 16'o016706);
`MEM('o016106, 16'o175602);
`MEM('o016110, 16'o104402);
`MEM('o016112, 16'o012767);
`MEM('o016114, 16'o016126);
`MEM('o016116, 16'o161664);
`MEM('o016120, 16'o016701);
`MEM('o016122, 16'o161424);
`MEM('o016124, 16'o000402);
`MEM('o016126, 16'o005267);
`MEM('o016130, 16'o001332);
`MEM('o016132, 16'o012767);
`MEM('o016134, 16'o016146);
`MEM('o016136, 16'o161644);
`MEM('o016140, 16'o024646);
`MEM('o016142, 16'o012701);
`MEM('o016144, 16'o160000);
`MEM('o016146, 16'o022626);
`MEM('o016150, 16'o014111);
`MEM('o016152, 16'o162701);
`MEM('o016154, 16'o000302);
`MEM('o016156, 16'o010167);
`MEM('o016160, 16'o001300);
`MEM('o016162, 16'o012700);
`MEM('o016164, 16'o013540);
`MEM('o016166, 16'o104552);
`MEM('o016170, 16'o122702);
`MEM('o016172, 16'o000114);
`MEM('o016174, 16'o001433);
`MEM('o016176, 16'o122702);
`MEM('o016200, 16'o000104);
`MEM('o016202, 16'o001435);
`MEM('o016204, 16'o122702);
`MEM('o016206, 16'o000105);
`MEM('o016210, 16'o001430);
`MEM('o016212, 16'o122702);
`MEM('o016214, 16'o000110);
`MEM('o016216, 16'o001432);
`MEM('o016220, 16'o122702);
`MEM('o016222, 16'o000012);
`MEM('o016224, 16'o001503);
`MEM('o016226, 16'o104470);
`MEM('o016230, 16'o001030);
`MEM('o016232, 16'o005301);
`MEM('o016234, 16'o104410);
`MEM('o016236, 16'o010067);
`MEM('o016240, 16'o001206);
`MEM('o016242, 16'o104472);
`MEM('o016244, 16'o122702);
`MEM('o016246, 16'o000012);
`MEM('o016250, 16'o001471);
`MEM('o016252, 16'o122702);
`MEM('o016254, 16'o000054);
`MEM('o016256, 16'o001371);
`MEM('o016260, 16'o104472);
`MEM('o016262, 16'o000742);
`MEM('o016264, 16'o005267);
`MEM('o016266, 16'o001162);
`MEM('o016270, 16'o000764);
`MEM('o016272, 16'o005267);
`MEM('o016274, 16'o001160);
`MEM('o016276, 16'o005267);
`MEM('o016300, 16'o001152);
`MEM('o016302, 16'o000757);
`MEM('o016304, 16'o005367);
`MEM('o016306, 16'o001150);
`MEM('o016310, 16'o000754);
`MEM('o016312, 16'o005067);
`MEM('o016314, 16'o001132);
`MEM('o016316, 16'o005067);
`MEM('o016320, 16'o001130);
`MEM('o016322, 16'o005067);
`MEM('o016324, 16'o001126);
`MEM('o016326, 16'o005067);
`MEM('o016330, 16'o001124);
`MEM('o016332, 16'o005067);
`MEM('o016334, 16'o001122);
`MEM('o016336, 16'o012700);
`MEM('o016340, 16'o017304);
`MEM('o016342, 16'o104552);
`MEM('o016344, 16'o010367);
`MEM('o016346, 16'o001104);
`MEM('o016350, 16'o003405);
`MEM('o016352, 16'o012700);
`MEM('o016354, 16'o017234);
`MEM('o016356, 16'o104552);
`MEM('o016360, 16'o010367);
`MEM('o016362, 16'o001072);
`MEM('o016364, 16'o005767);
`MEM('o016366, 16'o001074);
`MEM('o016370, 16'o001005);
`MEM('o016372, 16'o012700);
`MEM('o016374, 16'o017350);
`MEM('o016376, 16'o104552);
`MEM('o016400, 16'o010367);
`MEM('o016402, 16'o001046);
`MEM('o016404, 16'o012700);
`MEM('o016406, 16'o017401);
`MEM('o016410, 16'o104552);
`MEM('o016412, 16'o010367);
`MEM('o016414, 16'o001042);
`MEM('o016416, 16'o012700);
`MEM('o016420, 16'o017437);
`MEM('o016422, 16'o104466);
`MEM('o016424, 16'o104500);
`MEM('o016426, 16'o104410);
`MEM('o016430, 16'o010067);
`MEM('o016432, 16'o001014);
`MEM('o016434, 16'o066767);
`MEM('o016436, 16'o001024);
`MEM('o016440, 16'o001010);
`MEM('o016442, 16'o005767);
`MEM('o016444, 16'o001004);
`MEM('o016446, 16'o003407);
`MEM('o016450, 16'o012767);
`MEM('o016452, 16'o177560);
`MEM('o016454, 16'o175226);
`MEM('o016456, 16'o012767);
`MEM('o016460, 16'o177564);
`MEM('o016462, 16'o175222);
`MEM('o016464, 16'o000406);
`MEM('o016466, 16'o012767);
`MEM('o016470, 16'o177550);
`MEM('o016472, 16'o175210);
`MEM('o016474, 16'o012767);
`MEM('o016476, 16'o177554);
`MEM('o016500, 16'o175204);
`MEM('o016502, 16'o016701);
`MEM('o016504, 16'o000754);
`MEM('o016506, 16'o016700);
`MEM('o016510, 16'o000736);
`MEM('o016512, 16'o001414);
`MEM('o016514, 16'o000300);
`MEM('o016516, 16'o006300);
`MEM('o016520, 16'o006300);
`MEM('o016522, 16'o006300);
`MEM('o016524, 16'o042700);
`MEM('o016526, 16'o003777);
`MEM('o016530, 16'o020027);
`MEM('o016532, 16'o020000);
`MEM('o016534, 16'o103666);
`MEM('o016536, 16'o020001);
`MEM('o016540, 16'o101001);
`MEM('o016542, 16'o010001);
`MEM('o016544, 16'o010106);
`MEM('o016546, 16'o012767);
`MEM('o016550, 16'o000006);
`MEM('o016552, 16'o161230);
`MEM('o016554, 16'o010167);
`MEM('o016556, 16'o175132);
`MEM('o016560, 16'o012701);
`MEM('o016562, 16'o016104);
`MEM('o016564, 16'o005767);
`MEM('o016566, 16'o000664);
`MEM('o016570, 16'o003433);
`MEM('o016572, 16'o005067);
`MEM('o016574, 16'o167136);
`MEM('o016576, 16'o005067);
`MEM('o016600, 16'o167134);
`MEM('o016602, 16'o005067);
`MEM('o016604, 16'o167132);
`MEM('o016606, 16'o005067);
`MEM('o016610, 16'o167136);
`MEM('o016612, 16'o012701);
`MEM('o016614, 16'o015020);
`MEM('o016616, 16'o005767);
`MEM('o016620, 16'o000634);
`MEM('o016622, 16'o003416);
`MEM('o016624, 16'o005067);
`MEM('o016626, 16'o167112);
`MEM('o016630, 16'o005067);
`MEM('o016632, 16'o167110);
`MEM('o016634, 16'o012700);
`MEM('o016636, 16'o000136);
`MEM('o016640, 16'o006200);
`MEM('o016642, 16'o012701);
`MEM('o016644, 16'o013714);
`MEM('o016646, 16'o012702);
`MEM('o016650, 16'o017046);
`MEM('o016652, 16'o012221);
`MEM('o016654, 16'o005300);
`MEM('o016656, 16'o003375);
`MEM('o016660, 16'o005767);
`MEM('o016662, 16'o000574);
`MEM('o016664, 16'o002036);
`MEM('o016666, 16'o012767);
`MEM('o016670, 16'o016702);
`MEM('o016672, 16'o161160);
`MEM('o016674, 16'o010167);
`MEM('o016676, 16'o175002);
`MEM('o016700, 16'o000000);
`MEM('o016702, 16'o016701);
`MEM('o016704, 16'o174774);
`MEM('o016706, 16'o012700);
`MEM('o016710, 16'o000030);
`MEM('o016712, 16'o006200);
`MEM('o016714, 16'o012702);
`MEM('o016716, 16'o017204);
`MEM('o016720, 16'o010167);
`MEM('o016722, 16'o167062);
`MEM('o016724, 16'o010167);
`MEM('o016726, 16'o166514);
`MEM('o016730, 16'o012703);
`MEM('o016732, 16'o000016);
`MEM('o016734, 16'o060103);
`MEM('o016736, 16'o010367);
`MEM('o016740, 16'o161112);
`MEM('o016742, 16'o012221);
`MEM('o016744, 16'o005300);
`MEM('o016746, 16'o003375);
`MEM('o016750, 16'o016706);
`MEM('o016752, 16'o161074);
`MEM('o016754, 16'o010667);
`MEM('o016756, 16'o174732);
`MEM('o016760, 16'o000402);
`MEM('o016762, 16'o005067);
`MEM('o016764, 16'o166772);
`MEM('o016766, 16'o010167);
`MEM('o016770, 16'o174670);
`MEM('o016772, 16'o016705);
`MEM('o016774, 16'o174664);
`MEM('o016776, 16'o112725);
`MEM('o017000, 16'o000012);
`MEM('o017002, 16'o005067);
`MEM('o017004, 16'o174674);
`MEM('o017006, 16'o000167);
`MEM('o017010, 16'o164100);
`MEM('o017012, 16'o104466);
`MEM('o017014, 16'o104500);
`MEM('o017016, 16'o104472);
`MEM('o017020, 16'o005003);
`MEM('o017022, 16'o120227);
`MEM('o017024, 16'o000131);
`MEM('o017026, 16'o001002);
`MEM('o017030, 16'o005303);
`MEM('o017032, 16'o000207);
`MEM('o017034, 16'o120227);
`MEM('o017036, 16'o000116);
`MEM('o017040, 16'o001374);
`MEM('o017042, 16'o005203);
`MEM('o017044, 16'o000207);
`MEM('o017046, 16'o010046);
`MEM('o017050, 16'o104454);
`MEM('o017052, 16'o010100);
`MEM('o017054, 16'o104454);
`MEM('o017056, 16'o012701);
`MEM('o017060, 16'o010666);
`MEM('o017062, 16'o016600);
`MEM('o017064, 16'o000014);
`MEM('o017066, 16'o104432);
`MEM('o017070, 16'o010600);
`MEM('o017072, 16'o010046);
`MEM('o017074, 16'o010046);
`MEM('o017076, 16'o062716);
`MEM('o017100, 16'o000006);
`MEM('o017102, 16'o016600);
`MEM('o017104, 16'o000002);
`MEM('o017106, 16'o010001);
`MEM('o017110, 16'o004737);
`MEM('o017112, 16'o013372);
`MEM('o017114, 16'o005766);
`MEM('o017116, 16'o000006);
`MEM('o017120, 16'o003005);
`MEM('o017122, 16'o002416);
`MEM('o017124, 16'o062706);
`MEM('o017126, 16'o000022);
`MEM('o017130, 16'o000242);
`MEM('o017132, 16'o000207);
`MEM('o017134, 16'o011601);
`MEM('o017136, 16'o016600);
`MEM('o017140, 16'o000020);
`MEM('o017142, 16'o104430);
`MEM('o017144, 16'o012701);
`MEM('o017146, 16'o010666);
`MEM('o017150, 16'o016600);
`MEM('o017152, 16'o000002);
`MEM('o017154, 16'o104422);
`MEM('o017156, 16'o000756);
`MEM('o017160, 16'o011601);
`MEM('o017162, 16'o016600);
`MEM('o017164, 16'o000020);
`MEM('o017166, 16'o104426);
`MEM('o017170, 16'o012701);
`MEM('o017172, 16'o010666);
`MEM('o017174, 16'o016600);
`MEM('o017176, 16'o000002);
`MEM('o017200, 16'o104420);
`MEM('o017202, 16'o000744);
`MEM('o017204, 16'o062706);
`MEM('o017206, 16'o000010);
`MEM('o017210, 16'o010100);
`MEM('o017212, 16'o012601);
`MEM('o017214, 16'o013702);
`MEM('o017216, 16'o000050);
`MEM('o017220, 16'o000112);
`MEM('o017222, 16'o012602);
`MEM('o017224, 16'o012603);
`MEM('o017226, 16'o012604);
`MEM('o017230, 16'o000137);
`MEM('o017232, 16'o005430);
`MEM('o017234, 16'o047504);
`MEM('o017236, 16'o054440);
`MEM('o017240, 16'o052517);
`MEM('o017242, 16'o051040);
`MEM('o017244, 16'o050505);
`MEM('o017246, 16'o044525);
`MEM('o017250, 16'o042522);
`MEM('o017252, 16'o042440);
`MEM('o017254, 16'o050130);
`MEM('o017256, 16'o047440);
`MEM('o017260, 16'o020122);
`MEM('o017262, 16'o047514);
`MEM('o017264, 16'o020107);
`MEM('o017266, 16'o043050);
`MEM('o017270, 16'o047514);
`MEM('o017272, 16'o052101);
`MEM('o017274, 16'o047111);
`MEM('o017276, 16'o020107);
`MEM('o017300, 16'o024536);
`MEM('o017302, 16'o000077);
`MEM('o017304, 16'o047504);
`MEM('o017306, 16'o054440);
`MEM('o017310, 16'o052517);
`MEM('o017312, 16'o047040);
`MEM('o017314, 16'o042505);
`MEM('o017316, 16'o020104);
`MEM('o017320, 16'o044124);
`MEM('o017322, 16'o020105);
`MEM('o017324, 16'o054105);
`MEM('o017326, 16'o042524);
`MEM('o017330, 16'o042116);
`MEM('o017332, 16'o042105);
`MEM('o017334, 16'o043040);
`MEM('o017336, 16'o047125);
`MEM('o017340, 16'o052103);
`MEM('o017342, 16'o047511);
`MEM('o017344, 16'o051516);
`MEM('o017346, 16'o000077);
`MEM('o017350, 16'o044510);
`MEM('o017352, 16'o044107);
`MEM('o017354, 16'o051455);
`MEM('o017356, 16'o042520);
`MEM('o017360, 16'o042105);
`MEM('o017362, 16'o051040);
`MEM('o017364, 16'o040505);
`MEM('o017366, 16'o042504);
`MEM('o017370, 16'o027522);
`MEM('o017372, 16'o052520);
`MEM('o017374, 16'o041516);
`MEM('o017376, 16'o037510);
`MEM('o017400, 16'o051400);
`MEM('o017402, 16'o052105);
`MEM('o017404, 16'o052440);
`MEM('o017406, 16'o020120);
`MEM('o017410, 16'o044124);
`MEM('o017412, 16'o020105);
`MEM('o017414, 16'o054105);
`MEM('o017416, 16'o042524);
`MEM('o017420, 16'o047122);
`MEM('o017422, 16'o046101);
`MEM('o017424, 16'o043040);
`MEM('o017426, 16'o047125);
`MEM('o017430, 16'o052103);
`MEM('o017432, 16'o047511);
`MEM('o017434, 16'o037516);
`MEM('o017436, 16'o046400);
`MEM('o017440, 16'o046505);
`MEM('o017442, 16'o051117);
`MEM('o017444, 16'o037531);
`MEM('o017446, 16'o000000);
`MEM('o017450, 16'o000000);
`MEM('o017452, 16'o000000);
`MEM('o017454, 16'o000000);
`MEM('o017456, 16'o000000);
`MEM('o017460, 16'o000000);
`MEM('o017462, 16'o077474);
`MEM('o017464, 16'o000000);
`MEM('o017466, 16'o000000);
`MEM('o017470, 16'o000000);
`MEM('o017472, 16'o000000);
`MEM('o017474, 16'o000000);
`MEM('o017476, 16'o000000);
`MEM('o017500, 16'o000000);
`MEM('o017502, 16'o000000);
`MEM('o017504, 16'o000000);
`MEM('o017506, 16'o000000);
`MEM('o017510, 16'o000000);
`MEM('o017512, 16'o000000);
`MEM('o017514, 16'o000000);
`MEM('o017516, 16'o000000);
`MEM('o017520, 16'o000000);
`MEM('o017522, 16'o000000);
`MEM('o017524, 16'o000000);
`MEM('o017526, 16'o000000);
`MEM('o017530, 16'o000000);
`MEM('o017532, 16'o000000);
`MEM('o017534, 16'o000000);
`MEM('o017536, 16'o000000);
`MEM('o017540, 16'o000000);
`MEM('o017542, 16'o000000);
`MEM('o017544, 16'o000000);
`MEM('o017546, 16'o000000);
`MEM('o017550, 16'o000000);
`MEM('o017552, 16'o000000);
`MEM('o017554, 16'o000000);
`MEM('o017556, 16'o000000);
`MEM('o017560, 16'o000000);
`MEM('o017562, 16'o000000);
`MEM('o017564, 16'o000000);
`MEM('o017566, 16'o000000);
`MEM('o017570, 16'o000000);
`MEM('o017572, 16'o000000);
`MEM('o017574, 16'o000000);
`MEM('o017576, 16'o000000);
`MEM('o017600, 16'o000000);
`MEM('o017602, 16'o000000);
`MEM('o017604, 16'o000000);
`MEM('o017606, 16'o000000);
`MEM('o017610, 16'o000000);
`MEM('o017612, 16'o000000);
`MEM('o017614, 16'o000000);
`MEM('o017616, 16'o000000);
`MEM('o017620, 16'o000000);
`MEM('o017622, 16'o000000);
`MEM('o017624, 16'o000000);
`MEM('o017626, 16'o000000);
`MEM('o017630, 16'o000000);
`MEM('o017632, 16'o000000);
`MEM('o017634, 16'o000000);
`MEM('o017636, 16'o000000);
`MEM('o017640, 16'o000000);
`MEM('o017642, 16'o000000);
`MEM('o017644, 16'o000000);
`MEM('o017646, 16'o000000);
`MEM('o017650, 16'o000000);
`MEM('o017652, 16'o000000);
`MEM('o017654, 16'o000000);
`MEM('o017656, 16'o000000);
`MEM('o017660, 16'o000000);
`MEM('o017662, 16'o000000);
`MEM('o017664, 16'o000000);
`MEM('o017666, 16'o000000);
`MEM('o017670, 16'o000000);
`MEM('o017672, 16'o000000);
`MEM('o017674, 16'o000000);
`MEM('o017676, 16'o000000);
`MEM('o017700, 16'o000000);
`MEM('o017702, 16'o000000);
`MEM('o017704, 16'o000000);
`MEM('o017706, 16'o000000);
`MEM('o017710, 16'o000000);
`MEM('o017712, 16'o000000);
`MEM('o017714, 16'o000000);
`MEM('o017716, 16'o000000);
`MEM('o017720, 16'o000000);
`MEM('o017722, 16'o000000);
`MEM('o017724, 16'o000000);
`MEM('o017726, 16'o000000);
`MEM('o017730, 16'o000000);
`MEM('o017732, 16'o000000);
`MEM('o017734, 16'o000000);
`MEM('o017736, 16'o000000);
`MEM('o017740, 16'o000000);
`MEM('o017742, 16'o000000);
`MEM('o017744, 16'o000000);
`MEM('o017746, 16'o000000);
`MEM('o017750, 16'o000000);
`MEM('o017752, 16'o000000);
`MEM('o017754, 16'o000000);
`MEM('o017756, 16'o000000);
`MEM('o017760, 16'o000000);
`MEM('o017762, 16'o000000);
`MEM('o017764, 16'o000000);
`MEM('o017766, 16'o000000);
`MEM('o017770, 16'o000000);
`MEM('o017772, 16'o000000);
`MEM('o017774, 16'o000000);
`MEM('o017776, 16'o000000);
`MEM('o020000, 16'o000000);
`MEM('o020002, 16'o000000);
`MEM('o020004, 16'o000000);
`MEM('o020006, 16'o000000);
`MEM('o020010, 16'o000000);
`MEM('o020012, 16'o000000);
`MEM('o020014, 16'o000000);
`MEM('o020016, 16'o000000);
`MEM('o020020, 16'o000000);
`MEM('o020022, 16'o000000);
`MEM('o020024, 16'o000000);
`MEM('o020026, 16'o000000);
`MEM('o020030, 16'o000000);
`MEM('o020032, 16'o000000);
`MEM('o020034, 16'o000000);
`MEM('o020036, 16'o000000);
`MEM('o020040, 16'o000000);
`MEM('o020042, 16'o000000);
`MEM('o020044, 16'o000000);
`MEM('o020046, 16'o000000);
`MEM('o020050, 16'o000000);
`MEM('o020052, 16'o000000);
`MEM('o020054, 16'o000000);
`MEM('o020056, 16'o000000);
`MEM('o020060, 16'o000000);
`MEM('o020062, 16'o000000);
`MEM('o020064, 16'o000000);
`MEM('o020066, 16'o000000);
`MEM('o020070, 16'o000000);
`MEM('o020072, 16'o000000);
`MEM('o020074, 16'o000000);
`MEM('o020076, 16'o000000);
`MEM('o020100, 16'o000000);
`MEM('o020102, 16'o000000);
`MEM('o020104, 16'o000000);
`MEM('o020106, 16'o000000);
`MEM('o020110, 16'o000000);
`MEM('o020112, 16'o000000);
`MEM('o020114, 16'o000000);
`MEM('o020116, 16'o000000);
`MEM('o020120, 16'o000000);
`MEM('o020122, 16'o000000);
`MEM('o020124, 16'o000000);
`MEM('o020126, 16'o000000);
`MEM('o020130, 16'o000000);
`MEM('o020132, 16'o000000);
`MEM('o020134, 16'o000000);
`MEM('o020136, 16'o000000);
`MEM('o020140, 16'o000000);
`MEM('o020142, 16'o000000);
`MEM('o020144, 16'o000000);
`MEM('o020146, 16'o000000);
`MEM('o020150, 16'o000000);
`MEM('o020152, 16'o000000);
`MEM('o020154, 16'o000000);
`MEM('o020156, 16'o000000);
`MEM('o020160, 16'o000000);
`MEM('o020162, 16'o000000);
`MEM('o020164, 16'o000000);
`MEM('o020166, 16'o000000);
`MEM('o020170, 16'o000000);
`MEM('o020172, 16'o000000);
`MEM('o020174, 16'o000000);
`MEM('o020176, 16'o000000);
`MEM('o020200, 16'o000000);
`MEM('o020202, 16'o000000);
`MEM('o020204, 16'o000000);
`MEM('o020206, 16'o000000);
`MEM('o020210, 16'o000000);
`MEM('o020212, 16'o000000);
`MEM('o020214, 16'o000000);
`MEM('o020216, 16'o000000);
`MEM('o020220, 16'o000000);
`MEM('o020222, 16'o000000);
`MEM('o020224, 16'o000000);
`MEM('o020226, 16'o000000);
`MEM('o020230, 16'o000000);
`MEM('o020232, 16'o000000);
`MEM('o020234, 16'o000000);
`MEM('o020236, 16'o000000);
`MEM('o020240, 16'o000000);
`MEM('o020242, 16'o000000);
`MEM('o020244, 16'o000000);
`MEM('o020246, 16'o000000);
`MEM('o020250, 16'o000000);
`MEM('o020252, 16'o000000);
`MEM('o020254, 16'o000000);
`MEM('o020256, 16'o000000);
`MEM('o020260, 16'o000000);
`MEM('o020262, 16'o000000);
`MEM('o020264, 16'o000000);
`MEM('o020266, 16'o000000);
`MEM('o020270, 16'o000000);
`MEM('o020272, 16'o000000);
`MEM('o020274, 16'o000000);
`MEM('o020276, 16'o000000);
`MEM('o020300, 16'o000000);
`MEM('o020302, 16'o000000);
`MEM('o020304, 16'o000000);
`MEM('o020306, 16'o000000);
`MEM('o020310, 16'o000000);
`MEM('o020312, 16'o000000);
`MEM('o020314, 16'o000000);
`MEM('o020316, 16'o000000);
`MEM('o020320, 16'o000000);
`MEM('o020322, 16'o000000);
`MEM('o020324, 16'o000000);
`MEM('o020326, 16'o000000);
`MEM('o020330, 16'o000000);
`MEM('o020332, 16'o000000);
`MEM('o020334, 16'o000000);
`MEM('o020336, 16'o000000);
`MEM('o020340, 16'o000000);
`MEM('o020342, 16'o000000);
`MEM('o020344, 16'o000000);
`MEM('o020346, 16'o000000);
`MEM('o020350, 16'o000000);
`MEM('o020352, 16'o000000);
`MEM('o020354, 16'o000000);
`MEM('o020356, 16'o000000);
`MEM('o020360, 16'o000000);
`MEM('o020362, 16'o000000);
`MEM('o020364, 16'o000000);
`MEM('o020366, 16'o000000);
`MEM('o020370, 16'o000000);
`MEM('o020372, 16'o000000);
`MEM('o020374, 16'o000000);
`MEM('o020376, 16'o000000);
`MEM('o020400, 16'o000000);
`MEM('o020402, 16'o000000);
`MEM('o020404, 16'o000000);
`MEM('o020406, 16'o000000);
`MEM('o020410, 16'o000000);
`MEM('o020412, 16'o000000);
`MEM('o020414, 16'o000000);
`MEM('o020416, 16'o000000);
`MEM('o020420, 16'o000000);
`MEM('o020422, 16'o000000);
`MEM('o020424, 16'o000000);
`MEM('o020426, 16'o000000);
`MEM('o020430, 16'o000000);
`MEM('o020432, 16'o000000);
`MEM('o020434, 16'o000000);
`MEM('o020436, 16'o000000);
`MEM('o020440, 16'o000000);
`MEM('o020442, 16'o000000);
`MEM('o020444, 16'o000000);
`MEM('o020446, 16'o000000);
`MEM('o020450, 16'o000000);
`MEM('o020452, 16'o000000);
`MEM('o020454, 16'o000000);
`MEM('o020456, 16'o000000);
`MEM('o020460, 16'o000000);
`MEM('o020462, 16'o000000);
`MEM('o020464, 16'o000000);
`MEM('o020466, 16'o000000);
`MEM('o020470, 16'o000000);
`MEM('o020472, 16'o000000);
`MEM('o020474, 16'o000000);
`MEM('o020476, 16'o000000);
`MEM('o020500, 16'o000000);
`MEM('o020502, 16'o000000);
`MEM('o020504, 16'o000000);
`MEM('o020506, 16'o000000);
`MEM('o020510, 16'o000000);
`MEM('o020512, 16'o000000);
`MEM('o020514, 16'o000000);
`MEM('o020516, 16'o000000);
`MEM('o020520, 16'o000000);
`MEM('o020522, 16'o000000);
`MEM('o020524, 16'o000000);
`MEM('o020526, 16'o000000);
`MEM('o020530, 16'o000000);
`MEM('o020532, 16'o000000);
`MEM('o020534, 16'o000000);
`MEM('o020536, 16'o000000);
`MEM('o020540, 16'o000000);
`MEM('o020542, 16'o000000);
`MEM('o020544, 16'o000000);
`MEM('o020546, 16'o000000);
`MEM('o020550, 16'o000000);
`MEM('o020552, 16'o000000);
`MEM('o020554, 16'o000000);
`MEM('o020556, 16'o000000);
`MEM('o020560, 16'o000000);
`MEM('o020562, 16'o000000);
`MEM('o020564, 16'o000000);
`MEM('o020566, 16'o000000);
`MEM('o020570, 16'o000000);
`MEM('o020572, 16'o000000);
`MEM('o020574, 16'o000000);
`MEM('o020576, 16'o000000);
`MEM('o020600, 16'o000000);
`MEM('o020602, 16'o000000);
`MEM('o020604, 16'o000000);
`MEM('o020606, 16'o000000);
`MEM('o020610, 16'o000000);
`MEM('o020612, 16'o000000);
`MEM('o020614, 16'o000000);
`MEM('o020616, 16'o000000);
`MEM('o020620, 16'o000000);
`MEM('o020622, 16'o000000);
`MEM('o020624, 16'o000000);
`MEM('o020626, 16'o000000);
`MEM('o020630, 16'o000000);
`MEM('o020632, 16'o000000);
`MEM('o020634, 16'o000000);
`MEM('o020636, 16'o000000);
`MEM('o020640, 16'o000000);
`MEM('o020642, 16'o000000);
`MEM('o020644, 16'o000000);
`MEM('o020646, 16'o000000);
`MEM('o020650, 16'o000000);
`MEM('o020652, 16'o000000);
`MEM('o020654, 16'o000000);
`MEM('o020656, 16'o000000);
`MEM('o020660, 16'o000000);
`MEM('o020662, 16'o000000);
`MEM('o020664, 16'o000000);
`MEM('o020666, 16'o000000);
`MEM('o020670, 16'o000000);
`MEM('o020672, 16'o000000);
`MEM('o020674, 16'o000000);
`MEM('o020676, 16'o000000);
`MEM('o020700, 16'o000000);
`MEM('o020702, 16'o000000);
`MEM('o020704, 16'o000000);
`MEM('o020706, 16'o000000);
`MEM('o020710, 16'o000000);
`MEM('o020712, 16'o000000);
`MEM('o020714, 16'o000000);
`MEM('o020716, 16'o000000);
`MEM('o020720, 16'o000000);
`MEM('o020722, 16'o000000);
`MEM('o020724, 16'o000000);
`MEM('o020726, 16'o000000);
`MEM('o020730, 16'o000000);
`MEM('o020732, 16'o000000);
`MEM('o020734, 16'o000000);
`MEM('o020736, 16'o000000);
`MEM('o020740, 16'o000000);
`MEM('o020742, 16'o000000);
`MEM('o020744, 16'o000000);
`MEM('o020746, 16'o000000);
`MEM('o020750, 16'o000000);
`MEM('o020752, 16'o000000);
`MEM('o020754, 16'o000000);
`MEM('o020756, 16'o000000);
`MEM('o020760, 16'o000000);
`MEM('o020762, 16'o000000);
`MEM('o020764, 16'o000000);
`MEM('o020766, 16'o000000);
`MEM('o020770, 16'o000000);
`MEM('o020772, 16'o000000);
`MEM('o020774, 16'o000000);
`MEM('o020776, 16'o000000);
`MEM('o021000, 16'o000000);
`MEM('o021002, 16'o000000);
`MEM('o021004, 16'o000000);
`MEM('o021006, 16'o000000);
`MEM('o021010, 16'o000000);
`MEM('o021012, 16'o000000);
`MEM('o021014, 16'o000000);
`MEM('o021016, 16'o000000);
`MEM('o021020, 16'o000000);
`MEM('o021022, 16'o000000);
`MEM('o021024, 16'o000000);
`MEM('o021026, 16'o000000);
`MEM('o021030, 16'o000000);
`MEM('o021032, 16'o000000);
`MEM('o021034, 16'o000000);
`MEM('o021036, 16'o000000);
`MEM('o021040, 16'o000000);
`MEM('o021042, 16'o000000);
`MEM('o021044, 16'o000000);
`MEM('o021046, 16'o000000);
`MEM('o021050, 16'o000000);
`MEM('o021052, 16'o000000);
`MEM('o021054, 16'o000000);
`MEM('o021056, 16'o000000);
`MEM('o021060, 16'o000000);
`MEM('o021062, 16'o000000);
`MEM('o021064, 16'o000000);
`MEM('o021066, 16'o000000);
`MEM('o021070, 16'o000000);
`MEM('o021072, 16'o000000);
`MEM('o021074, 16'o000000);
`MEM('o021076, 16'o000000);
`MEM('o021100, 16'o000000);
`MEM('o021102, 16'o000000);
`MEM('o021104, 16'o000000);
`MEM('o021106, 16'o000000);
`MEM('o021110, 16'o000000);
`MEM('o021112, 16'o000000);
`MEM('o021114, 16'o000000);
`MEM('o021116, 16'o000000);
`MEM('o021120, 16'o000000);
`MEM('o021122, 16'o000000);
`MEM('o021124, 16'o000000);
`MEM('o021126, 16'o000000);
`MEM('o021130, 16'o000000);
`MEM('o021132, 16'o000000);
`MEM('o021134, 16'o000000);
`MEM('o021136, 16'o000000);
`MEM('o021140, 16'o000000);
`MEM('o021142, 16'o000000);
`MEM('o021144, 16'o000000);
`MEM('o021146, 16'o000000);
`MEM('o021150, 16'o000000);
`MEM('o021152, 16'o000000);
`MEM('o021154, 16'o000000);
`MEM('o021156, 16'o000000);
`MEM('o021160, 16'o000000);
`MEM('o021162, 16'o000000);
`MEM('o021164, 16'o000000);
`MEM('o021166, 16'o000000);
`MEM('o021170, 16'o000000);
`MEM('o021172, 16'o000000);
`MEM('o021174, 16'o000000);
`MEM('o021176, 16'o000000);
`MEM('o021200, 16'o000000);
`MEM('o021202, 16'o000000);
`MEM('o021204, 16'o000000);
`MEM('o021206, 16'o000000);
`MEM('o021210, 16'o000000);
`MEM('o021212, 16'o000000);
`MEM('o021214, 16'o000000);
`MEM('o021216, 16'o000000);
`MEM('o021220, 16'o000000);
`MEM('o021222, 16'o000000);
`MEM('o021224, 16'o000000);
`MEM('o021226, 16'o000000);
`MEM('o021230, 16'o000000);
`MEM('o021232, 16'o000000);
`MEM('o021234, 16'o000000);
`MEM('o021236, 16'o000000);
`MEM('o021240, 16'o000000);
`MEM('o021242, 16'o000000);
`MEM('o021244, 16'o000000);
`MEM('o021246, 16'o000000);
`MEM('o021250, 16'o000000);
`MEM('o021252, 16'o000000);
`MEM('o021254, 16'o000000);
`MEM('o021256, 16'o000000);
`MEM('o021260, 16'o000000);
`MEM('o021262, 16'o000000);
`MEM('o021264, 16'o000000);
`MEM('o021266, 16'o000000);
`MEM('o021270, 16'o000000);
`MEM('o021272, 16'o000000);
`MEM('o021274, 16'o000000);
`MEM('o021276, 16'o000000);
`MEM('o021300, 16'o000000);
`MEM('o021302, 16'o000000);
`MEM('o021304, 16'o000000);
`MEM('o021306, 16'o000000);
`MEM('o021310, 16'o000000);
`MEM('o021312, 16'o000000);
`MEM('o021314, 16'o000000);
`MEM('o021316, 16'o000000);
`MEM('o021320, 16'o000000);
`MEM('o021322, 16'o000000);
`MEM('o021324, 16'o000000);
`MEM('o021326, 16'o000000);
`MEM('o021330, 16'o000000);
`MEM('o021332, 16'o000000);
`MEM('o021334, 16'o000000);
`MEM('o021336, 16'o000000);
`MEM('o021340, 16'o000000);
`MEM('o021342, 16'o000000);
`MEM('o021344, 16'o000000);
`MEM('o021346, 16'o000000);
`MEM('o021350, 16'o000000);
`MEM('o021352, 16'o000000);
`MEM('o021354, 16'o000000);
`MEM('o021356, 16'o000000);
`MEM('o021360, 16'o000000);
`MEM('o021362, 16'o000000);
`MEM('o021364, 16'o000000);
`MEM('o021366, 16'o000000);
`MEM('o021370, 16'o000000);
`MEM('o021372, 16'o000000);
`MEM('o021374, 16'o000000);
`MEM('o021376, 16'o000000);
`MEM('o021400, 16'o000000);
`MEM('o021402, 16'o000000);
`MEM('o021404, 16'o000000);
`MEM('o021406, 16'o000000);
`MEM('o021410, 16'o000000);
`MEM('o021412, 16'o000000);
`MEM('o021414, 16'o000000);
`MEM('o021416, 16'o000000);
`MEM('o021420, 16'o000000);
`MEM('o021422, 16'o000000);
`MEM('o021424, 16'o000000);
`MEM('o021426, 16'o000000);
`MEM('o021430, 16'o000000);
`MEM('o021432, 16'o000000);
`MEM('o021434, 16'o000000);
`MEM('o021436, 16'o000000);
`MEM('o021440, 16'o000000);
`MEM('o021442, 16'o000000);
`MEM('o021444, 16'o000000);
`MEM('o021446, 16'o000000);
`MEM('o021450, 16'o000000);
`MEM('o021452, 16'o000000);
`MEM('o021454, 16'o000000);
`MEM('o021456, 16'o000000);
`MEM('o021460, 16'o000000);
`MEM('o021462, 16'o000000);
`MEM('o021464, 16'o000000);
`MEM('o021466, 16'o000000);
`MEM('o021470, 16'o000000);
`MEM('o021472, 16'o000000);
`MEM('o021474, 16'o000000);
`MEM('o021476, 16'o000000);
`MEM('o021500, 16'o000000);
`MEM('o021502, 16'o000000);
`MEM('o021504, 16'o000000);
`MEM('o021506, 16'o000000);
`MEM('o021510, 16'o000000);
`MEM('o021512, 16'o000000);
`MEM('o021514, 16'o000000);
`MEM('o021516, 16'o000000);
`MEM('o021520, 16'o000000);
`MEM('o021522, 16'o000000);
`MEM('o021524, 16'o000000);
`MEM('o021526, 16'o000000);
`MEM('o021530, 16'o000000);
`MEM('o021532, 16'o000000);
`MEM('o021534, 16'o000000);
`MEM('o021536, 16'o000000);
`MEM('o021540, 16'o000000);
`MEM('o021542, 16'o000000);
`MEM('o021544, 16'o000000);
`MEM('o021546, 16'o000000);
`MEM('o021550, 16'o000000);
`MEM('o021552, 16'o000000);
`MEM('o021554, 16'o000000);
`MEM('o021556, 16'o000000);
`MEM('o021560, 16'o000000);
`MEM('o021562, 16'o000000);
`MEM('o021564, 16'o000000);
`MEM('o021566, 16'o000000);
`MEM('o021570, 16'o000000);
`MEM('o021572, 16'o000000);
`MEM('o021574, 16'o000000);
`MEM('o021576, 16'o000000);
`MEM('o021600, 16'o000000);
`MEM('o021602, 16'o000000);
`MEM('o021604, 16'o000000);
`MEM('o021606, 16'o000000);
`MEM('o021610, 16'o000000);
`MEM('o021612, 16'o000000);
`MEM('o021614, 16'o000000);
`MEM('o021616, 16'o000000);
`MEM('o021620, 16'o000000);
`MEM('o021622, 16'o000000);
`MEM('o021624, 16'o000000);
`MEM('o021626, 16'o000000);
`MEM('o021630, 16'o000000);
`MEM('o021632, 16'o000000);
`MEM('o021634, 16'o000000);
`MEM('o021636, 16'o000000);
`MEM('o021640, 16'o000000);
`MEM('o021642, 16'o000000);
`MEM('o021644, 16'o000000);
`MEM('o021646, 16'o000000);
`MEM('o021650, 16'o000000);
`MEM('o021652, 16'o000000);
`MEM('o021654, 16'o000000);
`MEM('o021656, 16'o000000);
`MEM('o021660, 16'o000000);
`MEM('o021662, 16'o000000);
`MEM('o021664, 16'o000000);
`MEM('o021666, 16'o000000);
`MEM('o021670, 16'o000000);
`MEM('o021672, 16'o000000);
`MEM('o021674, 16'o000000);
`MEM('o021676, 16'o000000);
`MEM('o021700, 16'o000000);
`MEM('o021702, 16'o000000);
`MEM('o021704, 16'o000000);
`MEM('o021706, 16'o000000);
`MEM('o021710, 16'o000000);
`MEM('o021712, 16'o000000);
`MEM('o021714, 16'o000000);
`MEM('o021716, 16'o000000);
`MEM('o021720, 16'o000000);
`MEM('o021722, 16'o000000);
`MEM('o021724, 16'o000000);
`MEM('o021726, 16'o000000);
`MEM('o021730, 16'o000000);
`MEM('o021732, 16'o000000);
`MEM('o021734, 16'o000000);
`MEM('o021736, 16'o000000);
`MEM('o021740, 16'o000000);
`MEM('o021742, 16'o000000);
`MEM('o021744, 16'o000000);
`MEM('o021746, 16'o000000);
`MEM('o021750, 16'o000000);
`MEM('o021752, 16'o000000);
`MEM('o021754, 16'o000000);
`MEM('o021756, 16'o000000);
`MEM('o021760, 16'o000000);
`MEM('o021762, 16'o000000);
`MEM('o021764, 16'o000000);
`MEM('o021766, 16'o000000);
`MEM('o021770, 16'o000000);
`MEM('o021772, 16'o000000);
`MEM('o021774, 16'o000000);
`MEM('o021776, 16'o000000);
`MEM('o022000, 16'o000000);
`MEM('o022002, 16'o000000);
`MEM('o022004, 16'o000000);
`MEM('o022006, 16'o000000);
`MEM('o022010, 16'o000000);
`MEM('o022012, 16'o000000);
`MEM('o022014, 16'o000000);
`MEM('o022016, 16'o000000);
`MEM('o022020, 16'o000000);
`MEM('o022022, 16'o000000);
`MEM('o022024, 16'o000000);
`MEM('o022026, 16'o000000);
`MEM('o022030, 16'o000000);
`MEM('o022032, 16'o000000);
`MEM('o022034, 16'o000000);
`MEM('o022036, 16'o000000);
`MEM('o022040, 16'o000000);
`MEM('o022042, 16'o000000);
`MEM('o022044, 16'o000000);
`MEM('o022046, 16'o000000);
`MEM('o022050, 16'o000000);
`MEM('o022052, 16'o000000);
`MEM('o022054, 16'o000000);
`MEM('o022056, 16'o000000);
`MEM('o022060, 16'o000000);
`MEM('o022062, 16'o000000);
`MEM('o022064, 16'o000000);
`MEM('o022066, 16'o000000);
`MEM('o022070, 16'o000000);
`MEM('o022072, 16'o000000);
`MEM('o022074, 16'o000000);
`MEM('o022076, 16'o000000);
`MEM('o022100, 16'o000000);
`MEM('o022102, 16'o000000);
`MEM('o022104, 16'o000000);
`MEM('o022106, 16'o000000);
`MEM('o022110, 16'o000000);
`MEM('o022112, 16'o000000);
`MEM('o022114, 16'o000000);
`MEM('o022116, 16'o000000);
`MEM('o022120, 16'o000000);
`MEM('o022122, 16'o000000);
`MEM('o022124, 16'o000000);
`MEM('o022126, 16'o000000);
`MEM('o022130, 16'o000000);
`MEM('o022132, 16'o000000);
`MEM('o022134, 16'o000000);
`MEM('o022136, 16'o000000);
`MEM('o022140, 16'o000000);
`MEM('o022142, 16'o000000);
`MEM('o022144, 16'o000000);
`MEM('o022146, 16'o000000);
`MEM('o022150, 16'o000000);
`MEM('o022152, 16'o000000);
`MEM('o022154, 16'o000000);
`MEM('o022156, 16'o000000);
`MEM('o022160, 16'o000000);
`MEM('o022162, 16'o000000);
`MEM('o022164, 16'o000000);
`MEM('o022166, 16'o000000);
`MEM('o022170, 16'o000000);
`MEM('o022172, 16'o000000);
`MEM('o022174, 16'o000000);
`MEM('o022176, 16'o000000);
`MEM('o022200, 16'o000000);
`MEM('o022202, 16'o000000);
`MEM('o022204, 16'o000000);
`MEM('o022206, 16'o000000);
`MEM('o022210, 16'o000000);
`MEM('o022212, 16'o000000);
`MEM('o022214, 16'o000000);
`MEM('o022216, 16'o000000);
`MEM('o022220, 16'o000000);
`MEM('o022222, 16'o000000);
`MEM('o022224, 16'o000000);
`MEM('o022226, 16'o000000);
`MEM('o022230, 16'o000000);
`MEM('o022232, 16'o000000);
`MEM('o022234, 16'o000000);
`MEM('o022236, 16'o000000);
`MEM('o022240, 16'o000000);
`MEM('o022242, 16'o000000);
`MEM('o022244, 16'o000000);
`MEM('o022246, 16'o000000);
`MEM('o022250, 16'o000000);
`MEM('o022252, 16'o000000);
`MEM('o022254, 16'o000000);
`MEM('o022256, 16'o000000);
`MEM('o022260, 16'o000000);
`MEM('o022262, 16'o000000);
`MEM('o022264, 16'o000000);
`MEM('o022266, 16'o000000);
`MEM('o022270, 16'o000000);
`MEM('o022272, 16'o000000);
`MEM('o022274, 16'o000000);
`MEM('o022276, 16'o000000);
`MEM('o022300, 16'o000000);
`MEM('o022302, 16'o000000);
`MEM('o022304, 16'o000000);
`MEM('o022306, 16'o000000);
`MEM('o022310, 16'o000000);
`MEM('o022312, 16'o000000);
`MEM('o022314, 16'o000000);
`MEM('o022316, 16'o000000);
`MEM('o022320, 16'o000000);
`MEM('o022322, 16'o000000);
`MEM('o022324, 16'o000000);
`MEM('o022326, 16'o000000);
`MEM('o022330, 16'o000000);
`MEM('o022332, 16'o000000);
`MEM('o022334, 16'o000000);
`MEM('o022336, 16'o000000);
`MEM('o022340, 16'o000000);
`MEM('o022342, 16'o000000);
`MEM('o022344, 16'o000000);
`MEM('o022346, 16'o000000);
`MEM('o022350, 16'o000000);
`MEM('o022352, 16'o000000);
`MEM('o022354, 16'o000000);
`MEM('o022356, 16'o000000);
`MEM('o022360, 16'o000000);
`MEM('o022362, 16'o000000);
`MEM('o022364, 16'o000000);
`MEM('o022366, 16'o000000);
`MEM('o022370, 16'o000000);
`MEM('o022372, 16'o000000);
`MEM('o022374, 16'o000000);
`MEM('o022376, 16'o000000);
`MEM('o022400, 16'o000000);
`MEM('o022402, 16'o000000);
`MEM('o022404, 16'o000000);
`MEM('o022406, 16'o000000);
`MEM('o022410, 16'o000000);
`MEM('o022412, 16'o000000);
`MEM('o022414, 16'o000000);
`MEM('o022416, 16'o000000);
`MEM('o022420, 16'o000000);
`MEM('o022422, 16'o000000);
`MEM('o022424, 16'o000000);
`MEM('o022426, 16'o000000);
`MEM('o022430, 16'o000000);
`MEM('o022432, 16'o000000);
`MEM('o022434, 16'o000000);
`MEM('o022436, 16'o000000);
`MEM('o022440, 16'o000000);
`MEM('o022442, 16'o000000);
`MEM('o022444, 16'o000000);
`MEM('o022446, 16'o000000);
`MEM('o022450, 16'o000000);
`MEM('o022452, 16'o000000);
`MEM('o022454, 16'o000000);
`MEM('o022456, 16'o000000);
`MEM('o022460, 16'o000000);
`MEM('o022462, 16'o000000);
`MEM('o022464, 16'o000000);
`MEM('o022466, 16'o000000);
`MEM('o022470, 16'o000000);
`MEM('o022472, 16'o000000);
`MEM('o022474, 16'o000000);
`MEM('o022476, 16'o000000);
`MEM('o022500, 16'o000000);
`MEM('o022502, 16'o000000);
`MEM('o022504, 16'o000000);
`MEM('o022506, 16'o000000);
`MEM('o022510, 16'o000000);
`MEM('o022512, 16'o000000);
`MEM('o022514, 16'o000000);
`MEM('o022516, 16'o000000);
`MEM('o022520, 16'o000000);
`MEM('o022522, 16'o000000);
`MEM('o022524, 16'o000000);
`MEM('o022526, 16'o000000);
`MEM('o022530, 16'o000000);
`MEM('o022532, 16'o000000);
`MEM('o022534, 16'o000000);
`MEM('o022536, 16'o000000);
`MEM('o022540, 16'o000000);
`MEM('o022542, 16'o000000);
`MEM('o022544, 16'o000000);
`MEM('o022546, 16'o000000);
`MEM('o022550, 16'o000000);
`MEM('o022552, 16'o000000);
`MEM('o022554, 16'o000000);
`MEM('o022556, 16'o000000);
`MEM('o022560, 16'o000000);
`MEM('o022562, 16'o000000);
`MEM('o022564, 16'o000000);
`MEM('o022566, 16'o000000);
`MEM('o022570, 16'o000000);
`MEM('o022572, 16'o000000);
`MEM('o022574, 16'o000000);
`MEM('o022576, 16'o000000);
`MEM('o022600, 16'o000000);
`MEM('o022602, 16'o000000);
`MEM('o022604, 16'o000000);
`MEM('o022606, 16'o000000);
`MEM('o022610, 16'o000000);
`MEM('o022612, 16'o000000);
`MEM('o022614, 16'o000000);
`MEM('o022616, 16'o000000);
`MEM('o022620, 16'o000000);
`MEM('o022622, 16'o000000);
`MEM('o022624, 16'o000000);
`MEM('o022626, 16'o000000);
`MEM('o022630, 16'o000000);
`MEM('o022632, 16'o000000);
`MEM('o022634, 16'o000000);
`MEM('o022636, 16'o000000);
`MEM('o022640, 16'o000000);
`MEM('o022642, 16'o000000);
`MEM('o022644, 16'o000000);
`MEM('o022646, 16'o000000);
`MEM('o022650, 16'o000000);
`MEM('o022652, 16'o000000);
`MEM('o022654, 16'o000000);
`MEM('o022656, 16'o000000);
`MEM('o022660, 16'o000000);
`MEM('o022662, 16'o000000);
`MEM('o022664, 16'o000000);
`MEM('o022666, 16'o000000);
`MEM('o022670, 16'o000000);
`MEM('o022672, 16'o000000);
`MEM('o022674, 16'o000000);
`MEM('o022676, 16'o000000);
`MEM('o022700, 16'o000000);
`MEM('o022702, 16'o000000);
`MEM('o022704, 16'o000000);
`MEM('o022706, 16'o000000);
`MEM('o022710, 16'o000000);
`MEM('o022712, 16'o000000);
`MEM('o022714, 16'o000000);
`MEM('o022716, 16'o000000);
`MEM('o022720, 16'o000000);
`MEM('o022722, 16'o000000);
`MEM('o022724, 16'o000000);
`MEM('o022726, 16'o000000);
`MEM('o022730, 16'o000000);
`MEM('o022732, 16'o000000);
`MEM('o022734, 16'o000000);
`MEM('o022736, 16'o000000);
`MEM('o022740, 16'o000000);
`MEM('o022742, 16'o000000);
`MEM('o022744, 16'o000000);
`MEM('o022746, 16'o000000);
`MEM('o022750, 16'o000000);
`MEM('o022752, 16'o000000);
`MEM('o022754, 16'o000000);
`MEM('o022756, 16'o000000);
`MEM('o022760, 16'o000000);
`MEM('o022762, 16'o000000);
`MEM('o022764, 16'o000000);
`MEM('o022766, 16'o000000);
`MEM('o022770, 16'o000000);
`MEM('o022772, 16'o000000);
`MEM('o022774, 16'o000000);
`MEM('o022776, 16'o000000);
`MEM('o023000, 16'o000000);
`MEM('o023002, 16'o000000);
`MEM('o023004, 16'o000000);
`MEM('o023006, 16'o000000);
`MEM('o023010, 16'o000000);
`MEM('o023012, 16'o000000);
`MEM('o023014, 16'o000000);
`MEM('o023016, 16'o000000);
`MEM('o023020, 16'o000000);
`MEM('o023022, 16'o000000);
`MEM('o023024, 16'o000000);
`MEM('o023026, 16'o000000);
`MEM('o023030, 16'o000000);
`MEM('o023032, 16'o000000);
`MEM('o023034, 16'o000000);
`MEM('o023036, 16'o000000);
`MEM('o023040, 16'o000000);
`MEM('o023042, 16'o000000);
`MEM('o023044, 16'o000000);
`MEM('o023046, 16'o000000);
`MEM('o023050, 16'o000000);
`MEM('o023052, 16'o000000);
`MEM('o023054, 16'o000000);
`MEM('o023056, 16'o000000);
`MEM('o023060, 16'o000000);
`MEM('o023062, 16'o000000);
`MEM('o023064, 16'o000000);
`MEM('o023066, 16'o000000);
`MEM('o023070, 16'o000000);
`MEM('o023072, 16'o000000);
`MEM('o023074, 16'o000000);
`MEM('o023076, 16'o000000);
`MEM('o023100, 16'o000000);
`MEM('o023102, 16'o000000);
`MEM('o023104, 16'o000000);
`MEM('o023106, 16'o000000);
`MEM('o023110, 16'o000000);
`MEM('o023112, 16'o000000);
`MEM('o023114, 16'o000000);
`MEM('o023116, 16'o000000);
`MEM('o023120, 16'o000000);
`MEM('o023122, 16'o000000);
`MEM('o023124, 16'o000000);
`MEM('o023126, 16'o000000);
`MEM('o023130, 16'o000000);
`MEM('o023132, 16'o000000);
`MEM('o023134, 16'o000000);
`MEM('o023136, 16'o000000);
`MEM('o023140, 16'o000000);
`MEM('o023142, 16'o000000);
`MEM('o023144, 16'o000000);
`MEM('o023146, 16'o000000);
`MEM('o023150, 16'o000000);
`MEM('o023152, 16'o000000);
`MEM('o023154, 16'o000000);
`MEM('o023156, 16'o000000);
`MEM('o023160, 16'o000000);
`MEM('o023162, 16'o000000);
`MEM('o023164, 16'o000000);
`MEM('o023166, 16'o000000);
`MEM('o023170, 16'o000000);
`MEM('o023172, 16'o000000);
`MEM('o023174, 16'o000000);
`MEM('o023176, 16'o000000);
`MEM('o023200, 16'o000000);
`MEM('o023202, 16'o000000);
`MEM('o023204, 16'o000000);
`MEM('o023206, 16'o000000);
`MEM('o023210, 16'o000000);
`MEM('o023212, 16'o000000);
`MEM('o023214, 16'o000000);
`MEM('o023216, 16'o000000);
`MEM('o023220, 16'o000000);
`MEM('o023222, 16'o000000);
`MEM('o023224, 16'o000000);
`MEM('o023226, 16'o000000);
`MEM('o023230, 16'o000000);
`MEM('o023232, 16'o000000);
`MEM('o023234, 16'o000000);
`MEM('o023236, 16'o000000);
`MEM('o023240, 16'o000000);
`MEM('o023242, 16'o000000);
`MEM('o023244, 16'o000000);
`MEM('o023246, 16'o000000);
`MEM('o023250, 16'o000000);
`MEM('o023252, 16'o000000);
`MEM('o023254, 16'o000000);
`MEM('o023256, 16'o000000);
`MEM('o023260, 16'o000000);
`MEM('o023262, 16'o000000);
`MEM('o023264, 16'o000000);
`MEM('o023266, 16'o000000);
`MEM('o023270, 16'o000000);
`MEM('o023272, 16'o000000);
`MEM('o023274, 16'o000000);
`MEM('o023276, 16'o000000);
`MEM('o023300, 16'o000000);
`MEM('o023302, 16'o000000);
`MEM('o023304, 16'o000000);
`MEM('o023306, 16'o000000);
`MEM('o023310, 16'o000000);
`MEM('o023312, 16'o000000);
`MEM('o023314, 16'o000000);
`MEM('o023316, 16'o000000);
`MEM('o023320, 16'o000000);
`MEM('o023322, 16'o000000);
`MEM('o023324, 16'o000000);
`MEM('o023326, 16'o000000);
`MEM('o023330, 16'o000000);
`MEM('o023332, 16'o000000);
`MEM('o023334, 16'o000000);
`MEM('o023336, 16'o000000);
`MEM('o023340, 16'o000000);
`MEM('o023342, 16'o000000);
`MEM('o023344, 16'o000000);
`MEM('o023346, 16'o000000);
`MEM('o023350, 16'o000000);
`MEM('o023352, 16'o000000);
`MEM('o023354, 16'o000000);
`MEM('o023356, 16'o000000);
`MEM('o023360, 16'o000000);
`MEM('o023362, 16'o000000);
`MEM('o023364, 16'o000000);
`MEM('o023366, 16'o000000);
`MEM('o023370, 16'o000000);
`MEM('o023372, 16'o000000);
`MEM('o023374, 16'o000000);
`MEM('o023376, 16'o000000);
`MEM('o023400, 16'o000000);
`MEM('o023402, 16'o000000);
`MEM('o023404, 16'o000000);
`MEM('o023406, 16'o000000);
`MEM('o023410, 16'o000000);
`MEM('o023412, 16'o000000);
`MEM('o023414, 16'o000000);
`MEM('o023416, 16'o000000);
`MEM('o023420, 16'o000000);
`MEM('o023422, 16'o000000);
`MEM('o023424, 16'o000000);
`MEM('o023426, 16'o000000);
`MEM('o023430, 16'o000000);
`MEM('o023432, 16'o000000);
`MEM('o023434, 16'o000000);
`MEM('o023436, 16'o000000);
`MEM('o023440, 16'o000000);
`MEM('o023442, 16'o000000);
`MEM('o023444, 16'o000000);
`MEM('o023446, 16'o000000);
`MEM('o023450, 16'o000000);
`MEM('o023452, 16'o000000);
`MEM('o023454, 16'o000000);
`MEM('o023456, 16'o000000);
`MEM('o023460, 16'o000000);
`MEM('o023462, 16'o000000);
`MEM('o023464, 16'o000000);
`MEM('o023466, 16'o000000);
`MEM('o023470, 16'o000000);
`MEM('o023472, 16'o000000);
`MEM('o023474, 16'o000000);
`MEM('o023476, 16'o000000);
`MEM('o023500, 16'o000000);
`MEM('o023502, 16'o000000);
`MEM('o023504, 16'o000000);
`MEM('o023506, 16'o000000);
`MEM('o023510, 16'o000000);
`MEM('o023512, 16'o000000);
`MEM('o023514, 16'o000000);
`MEM('o023516, 16'o000000);
`MEM('o023520, 16'o000000);
`MEM('o023522, 16'o000000);
`MEM('o023524, 16'o000000);
`MEM('o023526, 16'o000000);
`MEM('o023530, 16'o000000);
`MEM('o023532, 16'o000000);
`MEM('o023534, 16'o000000);
`MEM('o023536, 16'o000000);
`MEM('o023540, 16'o000000);
`MEM('o023542, 16'o000000);
`MEM('o023544, 16'o000000);
`MEM('o023546, 16'o000000);
`MEM('o023550, 16'o000000);
`MEM('o023552, 16'o000000);
`MEM('o023554, 16'o000000);
`MEM('o023556, 16'o000000);
`MEM('o023560, 16'o000000);
`MEM('o023562, 16'o000000);
`MEM('o023564, 16'o000000);
`MEM('o023566, 16'o000000);
`MEM('o023570, 16'o000000);
`MEM('o023572, 16'o000000);
`MEM('o023574, 16'o000000);
`MEM('o023576, 16'o000000);
`MEM('o023600, 16'o000000);
`MEM('o023602, 16'o000000);
`MEM('o023604, 16'o000000);
`MEM('o023606, 16'o000000);
`MEM('o023610, 16'o000000);
`MEM('o023612, 16'o000000);
`MEM('o023614, 16'o000000);
`MEM('o023616, 16'o000000);
`MEM('o023620, 16'o000000);
`MEM('o023622, 16'o000000);
`MEM('o023624, 16'o000000);
`MEM('o023626, 16'o000000);
`MEM('o023630, 16'o000000);
`MEM('o023632, 16'o000000);
`MEM('o023634, 16'o000000);
`MEM('o023636, 16'o000000);
`MEM('o023640, 16'o000000);
`MEM('o023642, 16'o000000);
`MEM('o023644, 16'o000000);
`MEM('o023646, 16'o000000);
`MEM('o023650, 16'o000000);
`MEM('o023652, 16'o000000);
`MEM('o023654, 16'o000000);
`MEM('o023656, 16'o000000);
`MEM('o023660, 16'o000000);
`MEM('o023662, 16'o000000);
`MEM('o023664, 16'o000000);
`MEM('o023666, 16'o000000);
`MEM('o023670, 16'o000000);
`MEM('o023672, 16'o000000);
`MEM('o023674, 16'o000000);
`MEM('o023676, 16'o000000);
`MEM('o023700, 16'o000000);
`MEM('o023702, 16'o000000);
`MEM('o023704, 16'o000000);
`MEM('o023706, 16'o000000);
`MEM('o023710, 16'o000000);
`MEM('o023712, 16'o000000);
`MEM('o023714, 16'o000000);
`MEM('o023716, 16'o000000);
`MEM('o023720, 16'o000000);
`MEM('o023722, 16'o000000);
`MEM('o023724, 16'o000000);
`MEM('o023726, 16'o000000);
`MEM('o023730, 16'o000000);
`MEM('o023732, 16'o000000);
`MEM('o023734, 16'o000000);
`MEM('o023736, 16'o000000);
`MEM('o023740, 16'o000000);
`MEM('o023742, 16'o000000);
`MEM('o023744, 16'o000000);
`MEM('o023746, 16'o000000);
`MEM('o023750, 16'o000000);
`MEM('o023752, 16'o000000);
`MEM('o023754, 16'o000000);
`MEM('o023756, 16'o000000);
`MEM('o023760, 16'o000000);
`MEM('o023762, 16'o000000);
`MEM('o023764, 16'o000000);
`MEM('o023766, 16'o000000);
`MEM('o023770, 16'o000000);
`MEM('o023772, 16'o000000);
`MEM('o023774, 16'o000000);
`MEM('o023776, 16'o000000);
`MEM('o024000, 16'o000000);
`MEM('o024002, 16'o000000);
`MEM('o024004, 16'o000000);
`MEM('o024006, 16'o000000);
`MEM('o024010, 16'o000000);
`MEM('o024012, 16'o000000);
`MEM('o024014, 16'o000000);
`MEM('o024016, 16'o000000);
`MEM('o024020, 16'o000000);
`MEM('o024022, 16'o000000);
`MEM('o024024, 16'o000000);
`MEM('o024026, 16'o000000);
`MEM('o024030, 16'o000000);
`MEM('o024032, 16'o000000);
`MEM('o024034, 16'o000000);
`MEM('o024036, 16'o000000);
`MEM('o024040, 16'o000000);
`MEM('o024042, 16'o000000);
`MEM('o024044, 16'o000000);
`MEM('o024046, 16'o000000);
`MEM('o024050, 16'o000000);
`MEM('o024052, 16'o000000);
`MEM('o024054, 16'o000000);
`MEM('o024056, 16'o000000);
`MEM('o024060, 16'o000000);
`MEM('o024062, 16'o000000);
`MEM('o024064, 16'o000000);
`MEM('o024066, 16'o000000);
`MEM('o024070, 16'o000000);
`MEM('o024072, 16'o000000);
`MEM('o024074, 16'o000000);
`MEM('o024076, 16'o000000);
`MEM('o024100, 16'o000000);
`MEM('o024102, 16'o000000);
`MEM('o024104, 16'o000000);
`MEM('o024106, 16'o000000);
`MEM('o024110, 16'o000000);
`MEM('o024112, 16'o000000);
`MEM('o024114, 16'o000000);
`MEM('o024116, 16'o000000);
`MEM('o024120, 16'o000000);
`MEM('o024122, 16'o000000);
`MEM('o024124, 16'o000000);
`MEM('o024126, 16'o000000);
`MEM('o024130, 16'o000000);
`MEM('o024132, 16'o000000);
`MEM('o024134, 16'o000000);
`MEM('o024136, 16'o000000);
`MEM('o024140, 16'o000000);
`MEM('o024142, 16'o000000);
`MEM('o024144, 16'o000000);
`MEM('o024146, 16'o000000);
`MEM('o024150, 16'o000000);
`MEM('o024152, 16'o000000);
`MEM('o024154, 16'o000000);
`MEM('o024156, 16'o000000);
`MEM('o024160, 16'o000000);
`MEM('o024162, 16'o000000);
`MEM('o024164, 16'o000000);
`MEM('o024166, 16'o000000);
`MEM('o024170, 16'o000000);
`MEM('o024172, 16'o000000);
`MEM('o024174, 16'o000000);
`MEM('o024176, 16'o000000);
`MEM('o024200, 16'o000000);
`MEM('o024202, 16'o000000);
`MEM('o024204, 16'o000000);
`MEM('o024206, 16'o000000);
`MEM('o024210, 16'o000000);
`MEM('o024212, 16'o000000);
`MEM('o024214, 16'o000000);
`MEM('o024216, 16'o000000);
`MEM('o024220, 16'o000000);
`MEM('o024222, 16'o000000);
`MEM('o024224, 16'o000000);
`MEM('o024226, 16'o000000);
`MEM('o024230, 16'o000000);
`MEM('o024232, 16'o000000);
`MEM('o024234, 16'o000000);
`MEM('o024236, 16'o000000);
`MEM('o024240, 16'o000000);
`MEM('o024242, 16'o000000);
`MEM('o024244, 16'o000000);
`MEM('o024246, 16'o000000);
`MEM('o024250, 16'o000000);
`MEM('o024252, 16'o000000);
`MEM('o024254, 16'o000000);
`MEM('o024256, 16'o000000);
`MEM('o024260, 16'o000000);
`MEM('o024262, 16'o000000);
`MEM('o024264, 16'o000000);
`MEM('o024266, 16'o000000);
`MEM('o024270, 16'o000000);
`MEM('o024272, 16'o000000);
`MEM('o024274, 16'o000000);
`MEM('o024276, 16'o000000);
`MEM('o024300, 16'o000000);
`MEM('o024302, 16'o000000);
`MEM('o024304, 16'o000000);
`MEM('o024306, 16'o000000);
`MEM('o024310, 16'o000000);
`MEM('o024312, 16'o000000);
`MEM('o024314, 16'o000000);
`MEM('o024316, 16'o000000);
`MEM('o024320, 16'o000000);
`MEM('o024322, 16'o000000);
`MEM('o024324, 16'o000000);
`MEM('o024326, 16'o000000);
`MEM('o024330, 16'o000000);
`MEM('o024332, 16'o000000);
`MEM('o024334, 16'o000000);
`MEM('o024336, 16'o000000);
`MEM('o024340, 16'o000000);
`MEM('o024342, 16'o000000);
`MEM('o024344, 16'o000000);
`MEM('o024346, 16'o000000);
`MEM('o024350, 16'o000000);
`MEM('o024352, 16'o000000);
`MEM('o024354, 16'o000000);
`MEM('o024356, 16'o000000);
`MEM('o024360, 16'o000000);
`MEM('o024362, 16'o000000);
`MEM('o024364, 16'o000000);
`MEM('o024366, 16'o000000);
`MEM('o024370, 16'o000000);
`MEM('o024372, 16'o000000);
`MEM('o024374, 16'o000000);
`MEM('o024376, 16'o000000);
`MEM('o024400, 16'o000000);
`MEM('o024402, 16'o000000);
`MEM('o024404, 16'o000000);
`MEM('o024406, 16'o000000);
`MEM('o024410, 16'o000000);
`MEM('o024412, 16'o000000);
`MEM('o024414, 16'o000000);
`MEM('o024416, 16'o000000);
`MEM('o024420, 16'o000000);
`MEM('o024422, 16'o000000);
`MEM('o024424, 16'o000000);
`MEM('o024426, 16'o000000);
`MEM('o024430, 16'o000000);
`MEM('o024432, 16'o000000);
`MEM('o024434, 16'o000000);
`MEM('o024436, 16'o000000);
`MEM('o024440, 16'o000000);
`MEM('o024442, 16'o000000);
`MEM('o024444, 16'o000000);
`MEM('o024446, 16'o000000);
`MEM('o024450, 16'o000000);
`MEM('o024452, 16'o000000);
`MEM('o024454, 16'o000000);
`MEM('o024456, 16'o000000);
`MEM('o024460, 16'o000000);
`MEM('o024462, 16'o000000);
`MEM('o024464, 16'o000000);
`MEM('o024466, 16'o000000);
`MEM('o024470, 16'o000000);
`MEM('o024472, 16'o000000);
`MEM('o024474, 16'o000000);
`MEM('o024476, 16'o000000);
`MEM('o024500, 16'o000000);
`MEM('o024502, 16'o000000);
`MEM('o024504, 16'o000000);
`MEM('o024506, 16'o000000);
`MEM('o024510, 16'o000000);
`MEM('o024512, 16'o000000);
`MEM('o024514, 16'o000000);
`MEM('o024516, 16'o000000);
`MEM('o024520, 16'o000000);
`MEM('o024522, 16'o000000);
`MEM('o024524, 16'o000000);
`MEM('o024526, 16'o000000);
`MEM('o024530, 16'o000000);
`MEM('o024532, 16'o000000);
`MEM('o024534, 16'o000000);
`MEM('o024536, 16'o000000);
`MEM('o024540, 16'o000000);
`MEM('o024542, 16'o000000);
`MEM('o024544, 16'o000000);
`MEM('o024546, 16'o000000);
`MEM('o024550, 16'o000000);
`MEM('o024552, 16'o000000);
`MEM('o024554, 16'o000000);
`MEM('o024556, 16'o000000);
`MEM('o024560, 16'o000000);
`MEM('o024562, 16'o000000);
`MEM('o024564, 16'o000000);
`MEM('o024566, 16'o000000);
`MEM('o024570, 16'o000000);
`MEM('o024572, 16'o000000);
`MEM('o024574, 16'o000000);
`MEM('o024576, 16'o000000);
`MEM('o024600, 16'o000000);
`MEM('o024602, 16'o000000);
`MEM('o024604, 16'o000000);
`MEM('o024606, 16'o000000);
`MEM('o024610, 16'o000000);
`MEM('o024612, 16'o000000);
`MEM('o024614, 16'o000000);
`MEM('o024616, 16'o000000);
`MEM('o024620, 16'o000000);
`MEM('o024622, 16'o000000);
`MEM('o024624, 16'o000000);
`MEM('o024626, 16'o000000);
`MEM('o024630, 16'o000000);
`MEM('o024632, 16'o000000);
`MEM('o024634, 16'o000000);
`MEM('o024636, 16'o000000);
`MEM('o024640, 16'o000000);
`MEM('o024642, 16'o000000);
`MEM('o024644, 16'o000000);
`MEM('o024646, 16'o000000);
`MEM('o024650, 16'o000000);
`MEM('o024652, 16'o000000);
`MEM('o024654, 16'o000000);
`MEM('o024656, 16'o000000);
`MEM('o024660, 16'o000000);
`MEM('o024662, 16'o000000);
`MEM('o024664, 16'o000000);
`MEM('o024666, 16'o000000);
`MEM('o024670, 16'o000000);
`MEM('o024672, 16'o000000);
`MEM('o024674, 16'o000000);
`MEM('o024676, 16'o000000);
`MEM('o024700, 16'o000000);
`MEM('o024702, 16'o000000);
`MEM('o024704, 16'o000000);
`MEM('o024706, 16'o000000);
`MEM('o024710, 16'o000000);
`MEM('o024712, 16'o000000);
`MEM('o024714, 16'o000000);
`MEM('o024716, 16'o000000);
`MEM('o024720, 16'o000000);
`MEM('o024722, 16'o000000);
`MEM('o024724, 16'o000000);
`MEM('o024726, 16'o000000);
`MEM('o024730, 16'o000000);
`MEM('o024732, 16'o000000);
`MEM('o024734, 16'o000000);
`MEM('o024736, 16'o000000);
`MEM('o024740, 16'o000000);
`MEM('o024742, 16'o000000);
`MEM('o024744, 16'o000000);
`MEM('o024746, 16'o000000);
`MEM('o024750, 16'o000000);
`MEM('o024752, 16'o000000);
`MEM('o024754, 16'o000000);
`MEM('o024756, 16'o000000);
`MEM('o024760, 16'o000000);
`MEM('o024762, 16'o000000);
`MEM('o024764, 16'o000000);
`MEM('o024766, 16'o000000);
`MEM('o024770, 16'o000000);
`MEM('o024772, 16'o000000);
`MEM('o024774, 16'o000000);
`MEM('o024776, 16'o000000);
`MEM('o025000, 16'o000000);
`MEM('o025002, 16'o000000);
`MEM('o025004, 16'o000000);
`MEM('o025006, 16'o000000);
`MEM('o025010, 16'o000000);
`MEM('o025012, 16'o000000);
`MEM('o025014, 16'o000000);
`MEM('o025016, 16'o000000);
`MEM('o025020, 16'o000000);
`MEM('o025022, 16'o000000);
`MEM('o025024, 16'o000000);
`MEM('o025026, 16'o000000);
`MEM('o025030, 16'o000000);
`MEM('o025032, 16'o000000);
`MEM('o025034, 16'o000000);
`MEM('o025036, 16'o000000);
`MEM('o025040, 16'o000000);
`MEM('o025042, 16'o000000);
`MEM('o025044, 16'o000000);
`MEM('o025046, 16'o000000);
`MEM('o025050, 16'o000000);
`MEM('o025052, 16'o000000);
`MEM('o025054, 16'o000000);
`MEM('o025056, 16'o000000);
`MEM('o025060, 16'o000000);
`MEM('o025062, 16'o000000);
`MEM('o025064, 16'o000000);
`MEM('o025066, 16'o000000);
`MEM('o025070, 16'o000000);
`MEM('o025072, 16'o000000);
`MEM('o025074, 16'o000000);
`MEM('o025076, 16'o000000);
`MEM('o025100, 16'o000000);
`MEM('o025102, 16'o000000);
`MEM('o025104, 16'o000000);
`MEM('o025106, 16'o000000);
`MEM('o025110, 16'o000000);
`MEM('o025112, 16'o000000);
`MEM('o025114, 16'o000000);
`MEM('o025116, 16'o000000);
`MEM('o025120, 16'o000000);
`MEM('o025122, 16'o000000);
`MEM('o025124, 16'o000000);
`MEM('o025126, 16'o000000);
`MEM('o025130, 16'o000000);
`MEM('o025132, 16'o000000);
`MEM('o025134, 16'o000000);
`MEM('o025136, 16'o000000);
`MEM('o025140, 16'o000000);
`MEM('o025142, 16'o000000);
`MEM('o025144, 16'o000000);
`MEM('o025146, 16'o000000);
`MEM('o025150, 16'o000000);
`MEM('o025152, 16'o000000);
`MEM('o025154, 16'o000000);
`MEM('o025156, 16'o000000);
`MEM('o025160, 16'o000000);
`MEM('o025162, 16'o000000);
`MEM('o025164, 16'o000000);
`MEM('o025166, 16'o000000);
`MEM('o025170, 16'o000000);
`MEM('o025172, 16'o000000);
`MEM('o025174, 16'o000000);
`MEM('o025176, 16'o000000);
`MEM('o025200, 16'o000000);
`MEM('o025202, 16'o000000);
`MEM('o025204, 16'o000000);
`MEM('o025206, 16'o000000);
`MEM('o025210, 16'o000000);
`MEM('o025212, 16'o000000);
`MEM('o025214, 16'o000000);
`MEM('o025216, 16'o000000);
`MEM('o025220, 16'o000000);
`MEM('o025222, 16'o000000);
`MEM('o025224, 16'o000000);
`MEM('o025226, 16'o000000);
`MEM('o025230, 16'o000000);
`MEM('o025232, 16'o000000);
`MEM('o025234, 16'o000000);
`MEM('o025236, 16'o000000);
`MEM('o025240, 16'o000000);
`MEM('o025242, 16'o000000);
`MEM('o025244, 16'o000000);
`MEM('o025246, 16'o000000);
`MEM('o025250, 16'o000000);
`MEM('o025252, 16'o000000);
`MEM('o025254, 16'o000000);
`MEM('o025256, 16'o000000);
`MEM('o025260, 16'o000000);
`MEM('o025262, 16'o000000);
`MEM('o025264, 16'o000000);
`MEM('o025266, 16'o000000);
`MEM('o025270, 16'o000000);
`MEM('o025272, 16'o000000);
`MEM('o025274, 16'o000000);
`MEM('o025276, 16'o000000);
`MEM('o025300, 16'o000000);
`MEM('o025302, 16'o000000);
`MEM('o025304, 16'o000000);
`MEM('o025306, 16'o000000);
`MEM('o025310, 16'o000000);
`MEM('o025312, 16'o000000);
`MEM('o025314, 16'o000000);
`MEM('o025316, 16'o000000);
`MEM('o025320, 16'o000000);
`MEM('o025322, 16'o000000);
`MEM('o025324, 16'o000000);
`MEM('o025326, 16'o000000);
`MEM('o025330, 16'o000000);
`MEM('o025332, 16'o000000);
`MEM('o025334, 16'o000000);
`MEM('o025336, 16'o000000);
`MEM('o025340, 16'o000000);
`MEM('o025342, 16'o000000);
`MEM('o025344, 16'o000000);
`MEM('o025346, 16'o000000);
`MEM('o025350, 16'o000000);
`MEM('o025352, 16'o000000);
`MEM('o025354, 16'o000000);
`MEM('o025356, 16'o000000);
`MEM('o025360, 16'o000000);
`MEM('o025362, 16'o000000);
`MEM('o025364, 16'o000000);
`MEM('o025366, 16'o000000);
`MEM('o025370, 16'o000000);
`MEM('o025372, 16'o000000);
`MEM('o025374, 16'o000000);
`MEM('o025376, 16'o000000);
`MEM('o025400, 16'o000000);
`MEM('o025402, 16'o000000);
`MEM('o025404, 16'o000000);
`MEM('o025406, 16'o000000);
`MEM('o025410, 16'o000000);
`MEM('o025412, 16'o000000);
`MEM('o025414, 16'o000000);
`MEM('o025416, 16'o000000);
`MEM('o025420, 16'o000000);
`MEM('o025422, 16'o000000);
`MEM('o025424, 16'o000000);
`MEM('o025426, 16'o000000);
`MEM('o025430, 16'o000000);
`MEM('o025432, 16'o000000);
`MEM('o025434, 16'o000000);
`MEM('o025436, 16'o000000);
`MEM('o025440, 16'o000000);
`MEM('o025442, 16'o000000);
`MEM('o025444, 16'o000000);
`MEM('o025446, 16'o000000);
`MEM('o025450, 16'o000000);
`MEM('o025452, 16'o000000);
`MEM('o025454, 16'o000000);
`MEM('o025456, 16'o000000);
`MEM('o025460, 16'o000000);
`MEM('o025462, 16'o000000);
`MEM('o025464, 16'o000000);
`MEM('o025466, 16'o000000);
`MEM('o025470, 16'o000000);
`MEM('o025472, 16'o000000);
`MEM('o025474, 16'o000000);
`MEM('o025476, 16'o000000);
`MEM('o025500, 16'o000000);
`MEM('o025502, 16'o000000);
`MEM('o025504, 16'o000000);
`MEM('o025506, 16'o000000);
`MEM('o025510, 16'o000000);
`MEM('o025512, 16'o000000);
`MEM('o025514, 16'o000000);
`MEM('o025516, 16'o000000);
`MEM('o025520, 16'o000000);
`MEM('o025522, 16'o000000);
`MEM('o025524, 16'o000000);
`MEM('o025526, 16'o000000);
`MEM('o025530, 16'o000000);
`MEM('o025532, 16'o000000);
`MEM('o025534, 16'o000000);
`MEM('o025536, 16'o000000);
`MEM('o025540, 16'o000000);
`MEM('o025542, 16'o000000);
`MEM('o025544, 16'o000000);
`MEM('o025546, 16'o000000);
`MEM('o025550, 16'o000000);
`MEM('o025552, 16'o000000);
`MEM('o025554, 16'o000000);
`MEM('o025556, 16'o000000);
`MEM('o025560, 16'o000000);
`MEM('o025562, 16'o000000);
`MEM('o025564, 16'o000000);
`MEM('o025566, 16'o000000);
`MEM('o025570, 16'o000000);
`MEM('o025572, 16'o000000);
`MEM('o025574, 16'o000000);
`MEM('o025576, 16'o000000);
`MEM('o025600, 16'o000000);
`MEM('o025602, 16'o000000);
`MEM('o025604, 16'o000000);
`MEM('o025606, 16'o000000);
`MEM('o025610, 16'o000000);
`MEM('o025612, 16'o000000);
`MEM('o025614, 16'o000000);
`MEM('o025616, 16'o000000);
`MEM('o025620, 16'o000000);
`MEM('o025622, 16'o000000);
`MEM('o025624, 16'o000000);
`MEM('o025626, 16'o000000);
`MEM('o025630, 16'o000000);
`MEM('o025632, 16'o000000);
`MEM('o025634, 16'o000000);
`MEM('o025636, 16'o000000);
`MEM('o025640, 16'o000000);
`MEM('o025642, 16'o000000);
`MEM('o025644, 16'o000000);
`MEM('o025646, 16'o000000);
`MEM('o025650, 16'o000000);
`MEM('o025652, 16'o000000);
`MEM('o025654, 16'o000000);
`MEM('o025656, 16'o000000);
`MEM('o025660, 16'o000000);
`MEM('o025662, 16'o000000);
`MEM('o025664, 16'o000000);
`MEM('o025666, 16'o000000);
`MEM('o025670, 16'o000000);
`MEM('o025672, 16'o000000);
`MEM('o025674, 16'o000000);
`MEM('o025676, 16'o000000);
`MEM('o025700, 16'o000000);
`MEM('o025702, 16'o000000);
`MEM('o025704, 16'o000000);
`MEM('o025706, 16'o000000);
`MEM('o025710, 16'o000000);
`MEM('o025712, 16'o000000);
`MEM('o025714, 16'o000000);
`MEM('o025716, 16'o000000);
`MEM('o025720, 16'o000000);
`MEM('o025722, 16'o000000);
`MEM('o025724, 16'o000000);
`MEM('o025726, 16'o000000);
`MEM('o025730, 16'o000000);
`MEM('o025732, 16'o000000);
`MEM('o025734, 16'o000000);
`MEM('o025736, 16'o000000);
`MEM('o025740, 16'o000000);
`MEM('o025742, 16'o000000);
`MEM('o025744, 16'o000000);
`MEM('o025746, 16'o000000);
`MEM('o025750, 16'o000000);
`MEM('o025752, 16'o000000);
`MEM('o025754, 16'o000000);
`MEM('o025756, 16'o000000);
`MEM('o025760, 16'o000000);
`MEM('o025762, 16'o000000);
`MEM('o025764, 16'o000000);
`MEM('o025766, 16'o000000);
`MEM('o025770, 16'o000000);
`MEM('o025772, 16'o000000);
`MEM('o025774, 16'o000000);
`MEM('o025776, 16'o000000);
`MEM('o026000, 16'o000000);
`MEM('o026002, 16'o000000);
`MEM('o026004, 16'o000000);
`MEM('o026006, 16'o000000);
`MEM('o026010, 16'o000000);
`MEM('o026012, 16'o000000);
`MEM('o026014, 16'o000000);
`MEM('o026016, 16'o000000);
`MEM('o026020, 16'o000000);
`MEM('o026022, 16'o000000);
`MEM('o026024, 16'o000000);
`MEM('o026026, 16'o000000);
`MEM('o026030, 16'o000000);
`MEM('o026032, 16'o000000);
`MEM('o026034, 16'o000000);
`MEM('o026036, 16'o000000);
`MEM('o026040, 16'o000000);
`MEM('o026042, 16'o000000);
`MEM('o026044, 16'o000000);
`MEM('o026046, 16'o000000);
`MEM('o026050, 16'o000000);
`MEM('o026052, 16'o000000);
`MEM('o026054, 16'o000000);
`MEM('o026056, 16'o000000);
`MEM('o026060, 16'o000000);
`MEM('o026062, 16'o000000);
`MEM('o026064, 16'o000000);
`MEM('o026066, 16'o000000);
`MEM('o026070, 16'o000000);
`MEM('o026072, 16'o000000);
`MEM('o026074, 16'o000000);
`MEM('o026076, 16'o000000);
`MEM('o026100, 16'o000000);
`MEM('o026102, 16'o000000);
`MEM('o026104, 16'o000000);
`MEM('o026106, 16'o000000);
`MEM('o026110, 16'o000000);
`MEM('o026112, 16'o000000);
`MEM('o026114, 16'o000000);
`MEM('o026116, 16'o000000);
`MEM('o026120, 16'o000000);
`MEM('o026122, 16'o000000);
`MEM('o026124, 16'o000000);
`MEM('o026126, 16'o000000);
`MEM('o026130, 16'o000000);
`MEM('o026132, 16'o000000);
`MEM('o026134, 16'o000000);
`MEM('o026136, 16'o000000);
`MEM('o026140, 16'o000000);
`MEM('o026142, 16'o000000);
`MEM('o026144, 16'o000000);
`MEM('o026146, 16'o000000);
`MEM('o026150, 16'o000000);
`MEM('o026152, 16'o000000);
`MEM('o026154, 16'o000000);
`MEM('o026156, 16'o000000);
`MEM('o026160, 16'o000000);
`MEM('o026162, 16'o000000);
`MEM('o026164, 16'o000000);
`MEM('o026166, 16'o000000);
`MEM('o026170, 16'o000000);
`MEM('o026172, 16'o000000);
`MEM('o026174, 16'o000000);
`MEM('o026176, 16'o000000);
`MEM('o026200, 16'o000000);
`MEM('o026202, 16'o000000);
`MEM('o026204, 16'o000000);
`MEM('o026206, 16'o000000);
`MEM('o026210, 16'o000000);
`MEM('o026212, 16'o000000);
`MEM('o026214, 16'o000000);
`MEM('o026216, 16'o000000);
`MEM('o026220, 16'o000000);
`MEM('o026222, 16'o000000);
`MEM('o026224, 16'o000000);
`MEM('o026226, 16'o000000);
`MEM('o026230, 16'o000000);
`MEM('o026232, 16'o000000);
`MEM('o026234, 16'o000000);
`MEM('o026236, 16'o000000);
`MEM('o026240, 16'o000000);
`MEM('o026242, 16'o000000);
`MEM('o026244, 16'o000000);
`MEM('o026246, 16'o000000);
`MEM('o026250, 16'o000000);
`MEM('o026252, 16'o000000);
`MEM('o026254, 16'o000000);
`MEM('o026256, 16'o000000);
`MEM('o026260, 16'o000000);
`MEM('o026262, 16'o000000);
`MEM('o026264, 16'o000000);
`MEM('o026266, 16'o000000);
`MEM('o026270, 16'o000000);
`MEM('o026272, 16'o000000);
`MEM('o026274, 16'o000000);
`MEM('o026276, 16'o000000);
`MEM('o026300, 16'o000000);
`MEM('o026302, 16'o000000);
`MEM('o026304, 16'o000000);
`MEM('o026306, 16'o000000);
`MEM('o026310, 16'o000000);
`MEM('o026312, 16'o000000);
`MEM('o026314, 16'o000000);
`MEM('o026316, 16'o000000);
`MEM('o026320, 16'o000000);
`MEM('o026322, 16'o000000);
`MEM('o026324, 16'o000000);
`MEM('o026326, 16'o000000);
`MEM('o026330, 16'o000000);
`MEM('o026332, 16'o000000);
`MEM('o026334, 16'o000000);
`MEM('o026336, 16'o000000);
`MEM('o026340, 16'o000000);
`MEM('o026342, 16'o000000);
`MEM('o026344, 16'o000000);
`MEM('o026346, 16'o000000);
`MEM('o026350, 16'o000000);
`MEM('o026352, 16'o000000);
`MEM('o026354, 16'o000000);
`MEM('o026356, 16'o000000);
`MEM('o026360, 16'o000000);
`MEM('o026362, 16'o000000);
`MEM('o026364, 16'o000000);
`MEM('o026366, 16'o000000);
`MEM('o026370, 16'o000000);
`MEM('o026372, 16'o000000);
`MEM('o026374, 16'o000000);
`MEM('o026376, 16'o000000);
`MEM('o026400, 16'o000000);
`MEM('o026402, 16'o000000);
`MEM('o026404, 16'o000000);
`MEM('o026406, 16'o000000);
`MEM('o026410, 16'o000000);
`MEM('o026412, 16'o000000);
`MEM('o026414, 16'o000000);
`MEM('o026416, 16'o000000);
`MEM('o026420, 16'o000000);
`MEM('o026422, 16'o000000);
`MEM('o026424, 16'o000000);
`MEM('o026426, 16'o000000);
`MEM('o026430, 16'o000000);
`MEM('o026432, 16'o000000);
`MEM('o026434, 16'o000000);
`MEM('o026436, 16'o000000);
`MEM('o026440, 16'o000000);
`MEM('o026442, 16'o000000);
`MEM('o026444, 16'o000000);
`MEM('o026446, 16'o000000);
`MEM('o026450, 16'o000000);
`MEM('o026452, 16'o000000);
`MEM('o026454, 16'o000000);
`MEM('o026456, 16'o000000);
`MEM('o026460, 16'o000000);
`MEM('o026462, 16'o000000);
`MEM('o026464, 16'o000000);
`MEM('o026466, 16'o000000);
`MEM('o026470, 16'o000000);
`MEM('o026472, 16'o000000);
`MEM('o026474, 16'o000000);
`MEM('o026476, 16'o000000);
`MEM('o026500, 16'o000000);
`MEM('o026502, 16'o000000);
`MEM('o026504, 16'o000000);
`MEM('o026506, 16'o000000);
`MEM('o026510, 16'o000000);
`MEM('o026512, 16'o000000);
`MEM('o026514, 16'o000000);
`MEM('o026516, 16'o000000);
`MEM('o026520, 16'o000000);
`MEM('o026522, 16'o000000);
`MEM('o026524, 16'o000000);
`MEM('o026526, 16'o000000);
`MEM('o026530, 16'o000000);
`MEM('o026532, 16'o000000);
`MEM('o026534, 16'o000000);
`MEM('o026536, 16'o000000);
`MEM('o026540, 16'o000000);
`MEM('o026542, 16'o000000);
`MEM('o026544, 16'o000000);
`MEM('o026546, 16'o000000);
`MEM('o026550, 16'o000000);
`MEM('o026552, 16'o000000);
`MEM('o026554, 16'o000000);
`MEM('o026556, 16'o000000);
`MEM('o026560, 16'o000000);
`MEM('o026562, 16'o000000);
`MEM('o026564, 16'o000000);
`MEM('o026566, 16'o000000);
`MEM('o026570, 16'o000000);
`MEM('o026572, 16'o000000);
`MEM('o026574, 16'o000000);
`MEM('o026576, 16'o000000);
`MEM('o026600, 16'o000000);
`MEM('o026602, 16'o000000);
`MEM('o026604, 16'o000000);
`MEM('o026606, 16'o000000);
`MEM('o026610, 16'o000000);
`MEM('o026612, 16'o000000);
`MEM('o026614, 16'o000000);
`MEM('o026616, 16'o000000);
`MEM('o026620, 16'o000000);
`MEM('o026622, 16'o000000);
`MEM('o026624, 16'o000000);
`MEM('o026626, 16'o000000);
`MEM('o026630, 16'o000000);
`MEM('o026632, 16'o000000);
`MEM('o026634, 16'o000000);
`MEM('o026636, 16'o000000);
`MEM('o026640, 16'o000000);
`MEM('o026642, 16'o000000);
`MEM('o026644, 16'o000000);
`MEM('o026646, 16'o000000);
`MEM('o026650, 16'o000000);
`MEM('o026652, 16'o000000);
`MEM('o026654, 16'o000000);
`MEM('o026656, 16'o000000);
`MEM('o026660, 16'o000000);
`MEM('o026662, 16'o000000);
`MEM('o026664, 16'o000000);
`MEM('o026666, 16'o000000);
`MEM('o026670, 16'o000000);
`MEM('o026672, 16'o000000);
`MEM('o026674, 16'o000000);
`MEM('o026676, 16'o000000);
`MEM('o026700, 16'o000000);
`MEM('o026702, 16'o000000);
`MEM('o026704, 16'o000000);
`MEM('o026706, 16'o000000);
`MEM('o026710, 16'o000000);
`MEM('o026712, 16'o000000);
`MEM('o026714, 16'o000000);
`MEM('o026716, 16'o000000);
`MEM('o026720, 16'o000000);
`MEM('o026722, 16'o000000);
`MEM('o026724, 16'o000000);
`MEM('o026726, 16'o000000);
`MEM('o026730, 16'o000000);
`MEM('o026732, 16'o000000);
`MEM('o026734, 16'o000000);
`MEM('o026736, 16'o000000);
`MEM('o026740, 16'o000000);
`MEM('o026742, 16'o000000);
`MEM('o026744, 16'o000000);
`MEM('o026746, 16'o000000);
`MEM('o026750, 16'o000000);
`MEM('o026752, 16'o000000);
`MEM('o026754, 16'o000000);
`MEM('o026756, 16'o000000);
`MEM('o026760, 16'o000000);
`MEM('o026762, 16'o000000);
`MEM('o026764, 16'o000000);
`MEM('o026766, 16'o000000);
`MEM('o026770, 16'o000000);
`MEM('o026772, 16'o000000);
`MEM('o026774, 16'o000000);
`MEM('o026776, 16'o000000);
`MEM('o027000, 16'o000000);
`MEM('o027002, 16'o000000);
`MEM('o027004, 16'o000000);
`MEM('o027006, 16'o000000);
`MEM('o027010, 16'o000000);
`MEM('o027012, 16'o000000);
`MEM('o027014, 16'o000000);
`MEM('o027016, 16'o000000);
`MEM('o027020, 16'o000000);
`MEM('o027022, 16'o000000);
`MEM('o027024, 16'o000000);
`MEM('o027026, 16'o000000);
`MEM('o027030, 16'o000000);
`MEM('o027032, 16'o000000);
`MEM('o027034, 16'o000000);
`MEM('o027036, 16'o000000);
`MEM('o027040, 16'o000000);
`MEM('o027042, 16'o000000);
`MEM('o027044, 16'o000000);
`MEM('o027046, 16'o000000);
`MEM('o027050, 16'o000000);
`MEM('o027052, 16'o000000);
`MEM('o027054, 16'o000000);
`MEM('o027056, 16'o000000);
`MEM('o027060, 16'o000000);
`MEM('o027062, 16'o000000);
`MEM('o027064, 16'o000000);
`MEM('o027066, 16'o000000);
`MEM('o027070, 16'o000000);
`MEM('o027072, 16'o000000);
`MEM('o027074, 16'o000000);
`MEM('o027076, 16'o000000);
`MEM('o027100, 16'o000000);
`MEM('o027102, 16'o000000);
`MEM('o027104, 16'o000000);
`MEM('o027106, 16'o000000);
`MEM('o027110, 16'o000000);
`MEM('o027112, 16'o000000);
`MEM('o027114, 16'o000000);
`MEM('o027116, 16'o000000);
`MEM('o027120, 16'o000000);
`MEM('o027122, 16'o000000);
`MEM('o027124, 16'o000000);
`MEM('o027126, 16'o000000);
`MEM('o027130, 16'o000000);
`MEM('o027132, 16'o000000);
`MEM('o027134, 16'o000000);
`MEM('o027136, 16'o000000);
`MEM('o027140, 16'o000000);
`MEM('o027142, 16'o000000);
`MEM('o027144, 16'o000000);
`MEM('o027146, 16'o000000);
`MEM('o027150, 16'o000000);
`MEM('o027152, 16'o000000);
`MEM('o027154, 16'o000000);
`MEM('o027156, 16'o000000);
`MEM('o027160, 16'o000000);
`MEM('o027162, 16'o000000);
`MEM('o027164, 16'o000000);
`MEM('o027166, 16'o000000);
`MEM('o027170, 16'o000000);
`MEM('o027172, 16'o000000);
`MEM('o027174, 16'o000000);
`MEM('o027176, 16'o000000);
`MEM('o027200, 16'o000000);
`MEM('o027202, 16'o000000);
`MEM('o027204, 16'o000000);
`MEM('o027206, 16'o000000);
`MEM('o027210, 16'o000000);
`MEM('o027212, 16'o000000);
`MEM('o027214, 16'o000000);
`MEM('o027216, 16'o000000);
`MEM('o027220, 16'o000000);
`MEM('o027222, 16'o000000);
`MEM('o027224, 16'o000000);
`MEM('o027226, 16'o000000);
`MEM('o027230, 16'o000000);
`MEM('o027232, 16'o000000);
`MEM('o027234, 16'o000000);
`MEM('o027236, 16'o000000);
`MEM('o027240, 16'o000000);
`MEM('o027242, 16'o000000);
`MEM('o027244, 16'o000000);
`MEM('o027246, 16'o000000);
`MEM('o027250, 16'o000000);
`MEM('o027252, 16'o000000);
`MEM('o027254, 16'o000000);
`MEM('o027256, 16'o000000);
`MEM('o027260, 16'o000000);
`MEM('o027262, 16'o000000);
`MEM('o027264, 16'o000000);
`MEM('o027266, 16'o000000);
`MEM('o027270, 16'o000000);
`MEM('o027272, 16'o000000);
`MEM('o027274, 16'o000000);
`MEM('o027276, 16'o000000);
`MEM('o027300, 16'o000000);
`MEM('o027302, 16'o000000);
`MEM('o027304, 16'o000000);
`MEM('o027306, 16'o000000);
`MEM('o027310, 16'o000000);
`MEM('o027312, 16'o000000);
`MEM('o027314, 16'o000000);
`MEM('o027316, 16'o000000);
`MEM('o027320, 16'o000000);
`MEM('o027322, 16'o000000);
`MEM('o027324, 16'o000000);
`MEM('o027326, 16'o000000);
`MEM('o027330, 16'o000000);
`MEM('o027332, 16'o000000);
`MEM('o027334, 16'o000000);
`MEM('o027336, 16'o000000);
`MEM('o027340, 16'o000000);
`MEM('o027342, 16'o000000);
`MEM('o027344, 16'o000000);
`MEM('o027346, 16'o000000);
`MEM('o027350, 16'o000000);
`MEM('o027352, 16'o000000);
`MEM('o027354, 16'o000000);
`MEM('o027356, 16'o000000);
`MEM('o027360, 16'o000000);
`MEM('o027362, 16'o000000);
`MEM('o027364, 16'o000000);
`MEM('o027366, 16'o000000);
`MEM('o027370, 16'o000000);
`MEM('o027372, 16'o000000);
`MEM('o027374, 16'o000000);
`MEM('o027376, 16'o000000);
`MEM('o027400, 16'o000000);
`MEM('o027402, 16'o000000);
`MEM('o027404, 16'o000000);
`MEM('o027406, 16'o000000);
`MEM('o027410, 16'o000000);
`MEM('o027412, 16'o000000);
`MEM('o027414, 16'o000000);
`MEM('o027416, 16'o000000);
`MEM('o027420, 16'o000000);
`MEM('o027422, 16'o000000);
`MEM('o027424, 16'o000000);
`MEM('o027426, 16'o000000);
`MEM('o027430, 16'o000000);
`MEM('o027432, 16'o000000);
`MEM('o027434, 16'o000000);
`MEM('o027436, 16'o000000);
`MEM('o027440, 16'o000000);
`MEM('o027442, 16'o000000);
`MEM('o027444, 16'o000000);
`MEM('o027446, 16'o000000);
`MEM('o027450, 16'o000000);
`MEM('o027452, 16'o000000);
`MEM('o027454, 16'o000000);
`MEM('o027456, 16'o000000);
`MEM('o027460, 16'o000000);
`MEM('o027462, 16'o000000);
`MEM('o027464, 16'o000000);
`MEM('o027466, 16'o000000);
`MEM('o027470, 16'o000000);
`MEM('o027472, 16'o000000);
`MEM('o027474, 16'o000000);
`MEM('o027476, 16'o000000);
`MEM('o027500, 16'o000000);
`MEM('o027502, 16'o000000);
`MEM('o027504, 16'o000000);
`MEM('o027506, 16'o000000);
`MEM('o027510, 16'o000000);
`MEM('o027512, 16'o000000);
`MEM('o027514, 16'o000000);
`MEM('o027516, 16'o000000);
`MEM('o027520, 16'o000000);
`MEM('o027522, 16'o000000);
`MEM('o027524, 16'o000000);
`MEM('o027526, 16'o000000);
`MEM('o027530, 16'o000000);
`MEM('o027532, 16'o000000);
`MEM('o027534, 16'o000000);
`MEM('o027536, 16'o000000);
`MEM('o027540, 16'o000000);
`MEM('o027542, 16'o000000);
`MEM('o027544, 16'o000000);
`MEM('o027546, 16'o000000);
`MEM('o027550, 16'o000000);
`MEM('o027552, 16'o000000);
`MEM('o027554, 16'o000000);
`MEM('o027556, 16'o000000);
`MEM('o027560, 16'o000000);
`MEM('o027562, 16'o000000);
`MEM('o027564, 16'o000000);
`MEM('o027566, 16'o000000);
`MEM('o027570, 16'o000000);
`MEM('o027572, 16'o000000);
`MEM('o027574, 16'o000000);
`MEM('o027576, 16'o000000);
`MEM('o027600, 16'o000000);
`MEM('o027602, 16'o000000);
`MEM('o027604, 16'o000000);
`MEM('o027606, 16'o000000);
`MEM('o027610, 16'o000000);
`MEM('o027612, 16'o000000);
`MEM('o027614, 16'o000000);
`MEM('o027616, 16'o000000);
`MEM('o027620, 16'o000000);
`MEM('o027622, 16'o000000);
`MEM('o027624, 16'o000000);
`MEM('o027626, 16'o000000);
`MEM('o027630, 16'o000000);
`MEM('o027632, 16'o000000);
`MEM('o027634, 16'o000000);
`MEM('o027636, 16'o000000);
`MEM('o027640, 16'o000000);
`MEM('o027642, 16'o000000);
`MEM('o027644, 16'o000000);
`MEM('o027646, 16'o000000);
`MEM('o027650, 16'o000000);
`MEM('o027652, 16'o000000);
`MEM('o027654, 16'o000000);
`MEM('o027656, 16'o000000);
`MEM('o027660, 16'o000000);
`MEM('o027662, 16'o000000);
`MEM('o027664, 16'o000000);
`MEM('o027666, 16'o000000);
`MEM('o027670, 16'o000000);
`MEM('o027672, 16'o000000);
`MEM('o027674, 16'o000000);
`MEM('o027676, 16'o000000);
`MEM('o027700, 16'o000000);
`MEM('o027702, 16'o000000);
`MEM('o027704, 16'o000000);
`MEM('o027706, 16'o000000);
`MEM('o027710, 16'o000000);
`MEM('o027712, 16'o000000);
`MEM('o027714, 16'o000000);
`MEM('o027716, 16'o000000);
`MEM('o027720, 16'o000000);
`MEM('o027722, 16'o000000);
`MEM('o027724, 16'o000000);
`MEM('o027726, 16'o000000);
`MEM('o027730, 16'o000000);
`MEM('o027732, 16'o000000);
`MEM('o027734, 16'o000000);
`MEM('o027736, 16'o000000);
`MEM('o027740, 16'o000000);
`MEM('o027742, 16'o000000);
`MEM('o027744, 16'o000000);
`MEM('o027746, 16'o000000);
`MEM('o027750, 16'o000000);
`MEM('o027752, 16'o000000);
`MEM('o027754, 16'o000000);
`MEM('o027756, 16'o000000);
`MEM('o027760, 16'o000000);
`MEM('o027762, 16'o000000);
`MEM('o027764, 16'o000000);
`MEM('o027766, 16'o000000);
`MEM('o027770, 16'o000000);
`MEM('o027772, 16'o000000);
`MEM('o027774, 16'o000000);
`MEM('o027776, 16'o000000);
`MEM('o030000, 16'o000000);
`MEM('o030002, 16'o000000);
`MEM('o030004, 16'o000000);
`MEM('o030006, 16'o000000);
`MEM('o030010, 16'o000000);
`MEM('o030012, 16'o000000);
`MEM('o030014, 16'o000000);
`MEM('o030016, 16'o000000);
`MEM('o030020, 16'o000000);
`MEM('o030022, 16'o000000);
`MEM('o030024, 16'o000000);
`MEM('o030026, 16'o000000);
`MEM('o030030, 16'o000000);
`MEM('o030032, 16'o000000);
`MEM('o030034, 16'o000000);
`MEM('o030036, 16'o000000);
`MEM('o030040, 16'o000000);
`MEM('o030042, 16'o000000);
`MEM('o030044, 16'o000000);
`MEM('o030046, 16'o000000);
`MEM('o030050, 16'o000000);
`MEM('o030052, 16'o000000);
`MEM('o030054, 16'o000000);
`MEM('o030056, 16'o000000);
`MEM('o030060, 16'o000000);
`MEM('o030062, 16'o000000);
`MEM('o030064, 16'o000000);
`MEM('o030066, 16'o000000);
`MEM('o030070, 16'o000000);
`MEM('o030072, 16'o000000);
`MEM('o030074, 16'o000000);
`MEM('o030076, 16'o000000);
`MEM('o030100, 16'o000000);
`MEM('o030102, 16'o000000);
`MEM('o030104, 16'o000000);
`MEM('o030106, 16'o000000);
`MEM('o030110, 16'o000000);
`MEM('o030112, 16'o000000);
`MEM('o030114, 16'o000000);
`MEM('o030116, 16'o000000);
`MEM('o030120, 16'o000000);
`MEM('o030122, 16'o000000);
`MEM('o030124, 16'o000000);
`MEM('o030126, 16'o000000);
`MEM('o030130, 16'o000000);
`MEM('o030132, 16'o000000);
`MEM('o030134, 16'o000000);
`MEM('o030136, 16'o000000);
`MEM('o030140, 16'o000000);
`MEM('o030142, 16'o000000);
`MEM('o030144, 16'o000000);
`MEM('o030146, 16'o000000);
`MEM('o030150, 16'o000000);
`MEM('o030152, 16'o000000);
`MEM('o030154, 16'o000000);
`MEM('o030156, 16'o000000);
`MEM('o030160, 16'o000000);
`MEM('o030162, 16'o000000);
`MEM('o030164, 16'o000000);
`MEM('o030166, 16'o000000);
`MEM('o030170, 16'o000000);
`MEM('o030172, 16'o000000);
`MEM('o030174, 16'o000000);
`MEM('o030176, 16'o000000);
`MEM('o030200, 16'o000000);
`MEM('o030202, 16'o000000);
`MEM('o030204, 16'o000000);
`MEM('o030206, 16'o000000);
`MEM('o030210, 16'o000000);
`MEM('o030212, 16'o000000);
`MEM('o030214, 16'o000000);
`MEM('o030216, 16'o000000);
`MEM('o030220, 16'o000000);
`MEM('o030222, 16'o000000);
`MEM('o030224, 16'o000000);
`MEM('o030226, 16'o000000);
`MEM('o030230, 16'o000000);
`MEM('o030232, 16'o000000);
`MEM('o030234, 16'o000000);
`MEM('o030236, 16'o000000);
`MEM('o030240, 16'o000000);
`MEM('o030242, 16'o000000);
`MEM('o030244, 16'o000000);
`MEM('o030246, 16'o000000);
`MEM('o030250, 16'o000000);
`MEM('o030252, 16'o000000);
`MEM('o030254, 16'o000000);
`MEM('o030256, 16'o000000);
`MEM('o030260, 16'o000000);
`MEM('o030262, 16'o000000);
`MEM('o030264, 16'o000000);
`MEM('o030266, 16'o000000);
`MEM('o030270, 16'o000000);
`MEM('o030272, 16'o000000);
`MEM('o030274, 16'o000000);
`MEM('o030276, 16'o000000);
`MEM('o030300, 16'o000000);
`MEM('o030302, 16'o000000);
`MEM('o030304, 16'o000000);
`MEM('o030306, 16'o000000);
`MEM('o030310, 16'o000000);
`MEM('o030312, 16'o000000);
`MEM('o030314, 16'o000000);
`MEM('o030316, 16'o000000);
`MEM('o030320, 16'o000000);
`MEM('o030322, 16'o000000);
`MEM('o030324, 16'o000000);
`MEM('o030326, 16'o000000);
`MEM('o030330, 16'o000000);
`MEM('o030332, 16'o000000);
`MEM('o030334, 16'o000000);
`MEM('o030336, 16'o000000);
`MEM('o030340, 16'o000000);
`MEM('o030342, 16'o000000);
`MEM('o030344, 16'o000000);
`MEM('o030346, 16'o000000);
`MEM('o030350, 16'o000000);
`MEM('o030352, 16'o000000);
`MEM('o030354, 16'o000000);
`MEM('o030356, 16'o000000);
`MEM('o030360, 16'o000000);
`MEM('o030362, 16'o000000);
`MEM('o030364, 16'o000000);
`MEM('o030366, 16'o000000);
`MEM('o030370, 16'o000000);
`MEM('o030372, 16'o000000);
`MEM('o030374, 16'o000000);
`MEM('o030376, 16'o000000);
`MEM('o030400, 16'o000000);
`MEM('o030402, 16'o000000);
`MEM('o030404, 16'o000000);
`MEM('o030406, 16'o000000);
`MEM('o030410, 16'o000000);
`MEM('o030412, 16'o000000);
`MEM('o030414, 16'o000000);
`MEM('o030416, 16'o000000);
`MEM('o030420, 16'o000000);
`MEM('o030422, 16'o000000);
`MEM('o030424, 16'o000000);
`MEM('o030426, 16'o000000);
`MEM('o030430, 16'o000000);
`MEM('o030432, 16'o000000);
`MEM('o030434, 16'o000000);
`MEM('o030436, 16'o000000);
`MEM('o030440, 16'o000000);
`MEM('o030442, 16'o000000);
`MEM('o030444, 16'o000000);
`MEM('o030446, 16'o000000);
`MEM('o030450, 16'o000000);
`MEM('o030452, 16'o000000);
`MEM('o030454, 16'o000000);
`MEM('o030456, 16'o000000);
`MEM('o030460, 16'o000000);
`MEM('o030462, 16'o000000);
`MEM('o030464, 16'o000000);
`MEM('o030466, 16'o000000);
`MEM('o030470, 16'o000000);
`MEM('o030472, 16'o000000);
`MEM('o030474, 16'o000000);
`MEM('o030476, 16'o000000);
`MEM('o030500, 16'o000000);
`MEM('o030502, 16'o000000);
`MEM('o030504, 16'o000000);
`MEM('o030506, 16'o000000);
`MEM('o030510, 16'o000000);
`MEM('o030512, 16'o000000);
`MEM('o030514, 16'o000000);
`MEM('o030516, 16'o000000);
`MEM('o030520, 16'o000000);
`MEM('o030522, 16'o000000);
`MEM('o030524, 16'o000000);
`MEM('o030526, 16'o000000);
`MEM('o030530, 16'o000000);
`MEM('o030532, 16'o000000);
`MEM('o030534, 16'o000000);
`MEM('o030536, 16'o000000);
`MEM('o030540, 16'o000000);
`MEM('o030542, 16'o000000);
`MEM('o030544, 16'o000000);
`MEM('o030546, 16'o000000);
`MEM('o030550, 16'o000000);
`MEM('o030552, 16'o000000);
`MEM('o030554, 16'o000000);
`MEM('o030556, 16'o000000);
`MEM('o030560, 16'o000000);
`MEM('o030562, 16'o000000);
`MEM('o030564, 16'o000000);
`MEM('o030566, 16'o000000);
`MEM('o030570, 16'o000000);
`MEM('o030572, 16'o000000);
`MEM('o030574, 16'o000000);
`MEM('o030576, 16'o000000);
`MEM('o030600, 16'o000000);
`MEM('o030602, 16'o000000);
`MEM('o030604, 16'o000000);
`MEM('o030606, 16'o000000);
`MEM('o030610, 16'o000000);
`MEM('o030612, 16'o000000);
`MEM('o030614, 16'o000000);
`MEM('o030616, 16'o000000);
`MEM('o030620, 16'o000000);
`MEM('o030622, 16'o000000);
`MEM('o030624, 16'o000000);
`MEM('o030626, 16'o000000);
`MEM('o030630, 16'o000000);
`MEM('o030632, 16'o000000);
`MEM('o030634, 16'o000000);
`MEM('o030636, 16'o000000);
`MEM('o030640, 16'o000000);
`MEM('o030642, 16'o000000);
`MEM('o030644, 16'o000000);
`MEM('o030646, 16'o000000);
`MEM('o030650, 16'o000000);
`MEM('o030652, 16'o000000);
`MEM('o030654, 16'o000000);
`MEM('o030656, 16'o000000);
`MEM('o030660, 16'o000000);
`MEM('o030662, 16'o000000);
`MEM('o030664, 16'o000000);
`MEM('o030666, 16'o000000);
`MEM('o030670, 16'o000000);
`MEM('o030672, 16'o000000);
`MEM('o030674, 16'o000000);
`MEM('o030676, 16'o000000);
`MEM('o030700, 16'o000000);
`MEM('o030702, 16'o000000);
`MEM('o030704, 16'o000000);
`MEM('o030706, 16'o000000);
`MEM('o030710, 16'o000000);
`MEM('o030712, 16'o000000);
`MEM('o030714, 16'o000000);
`MEM('o030716, 16'o000000);
`MEM('o030720, 16'o000000);
`MEM('o030722, 16'o000000);
`MEM('o030724, 16'o000000);
`MEM('o030726, 16'o000000);
`MEM('o030730, 16'o000000);
`MEM('o030732, 16'o000000);
`MEM('o030734, 16'o000000);
`MEM('o030736, 16'o000000);
`MEM('o030740, 16'o000000);
`MEM('o030742, 16'o000000);
`MEM('o030744, 16'o000000);
`MEM('o030746, 16'o000000);
`MEM('o030750, 16'o000000);
`MEM('o030752, 16'o000000);
`MEM('o030754, 16'o000000);
`MEM('o030756, 16'o000000);
`MEM('o030760, 16'o000000);
`MEM('o030762, 16'o000000);
`MEM('o030764, 16'o000000);
`MEM('o030766, 16'o000000);
`MEM('o030770, 16'o000000);
`MEM('o030772, 16'o000000);
`MEM('o030774, 16'o000000);
`MEM('o030776, 16'o000000);
`MEM('o031000, 16'o000000);
`MEM('o031002, 16'o000000);
`MEM('o031004, 16'o000000);
`MEM('o031006, 16'o000000);
`MEM('o031010, 16'o000000);
`MEM('o031012, 16'o000000);
`MEM('o031014, 16'o000000);
`MEM('o031016, 16'o000000);
`MEM('o031020, 16'o000000);
`MEM('o031022, 16'o000000);
`MEM('o031024, 16'o000000);
`MEM('o031026, 16'o000000);
`MEM('o031030, 16'o000000);
`MEM('o031032, 16'o000000);
`MEM('o031034, 16'o000000);
`MEM('o031036, 16'o000000);
`MEM('o031040, 16'o000000);
`MEM('o031042, 16'o000000);
`MEM('o031044, 16'o000000);
`MEM('o031046, 16'o000000);
`MEM('o031050, 16'o000000);
`MEM('o031052, 16'o000000);
`MEM('o031054, 16'o000000);
`MEM('o031056, 16'o000000);
`MEM('o031060, 16'o000000);
`MEM('o031062, 16'o000000);
`MEM('o031064, 16'o000000);
`MEM('o031066, 16'o000000);
`MEM('o031070, 16'o000000);
`MEM('o031072, 16'o000000);
`MEM('o031074, 16'o000000);
`MEM('o031076, 16'o000000);
`MEM('o031100, 16'o000000);
`MEM('o031102, 16'o000000);
`MEM('o031104, 16'o000000);
`MEM('o031106, 16'o000000);
`MEM('o031110, 16'o000000);
`MEM('o031112, 16'o000000);
`MEM('o031114, 16'o000000);
`MEM('o031116, 16'o000000);
`MEM('o031120, 16'o000000);
`MEM('o031122, 16'o000000);
`MEM('o031124, 16'o000000);
`MEM('o031126, 16'o000000);
`MEM('o031130, 16'o000000);
`MEM('o031132, 16'o000000);
`MEM('o031134, 16'o000000);
`MEM('o031136, 16'o000000);
`MEM('o031140, 16'o000000);
`MEM('o031142, 16'o000000);
`MEM('o031144, 16'o000000);
`MEM('o031146, 16'o000000);
`MEM('o031150, 16'o000000);
`MEM('o031152, 16'o000000);
`MEM('o031154, 16'o000000);
`MEM('o031156, 16'o000000);
`MEM('o031160, 16'o000000);
`MEM('o031162, 16'o000000);
`MEM('o031164, 16'o000000);
`MEM('o031166, 16'o000000);
`MEM('o031170, 16'o000000);
`MEM('o031172, 16'o000000);
`MEM('o031174, 16'o000000);
`MEM('o031176, 16'o000000);
`MEM('o031200, 16'o000000);
`MEM('o031202, 16'o000000);
`MEM('o031204, 16'o000000);
`MEM('o031206, 16'o000000);
`MEM('o031210, 16'o000000);
`MEM('o031212, 16'o000000);
`MEM('o031214, 16'o000000);
`MEM('o031216, 16'o000000);
`MEM('o031220, 16'o000000);
`MEM('o031222, 16'o000000);
`MEM('o031224, 16'o000000);
`MEM('o031226, 16'o000000);
`MEM('o031230, 16'o000000);
`MEM('o031232, 16'o000000);
`MEM('o031234, 16'o000000);
`MEM('o031236, 16'o000000);
`MEM('o031240, 16'o000000);
`MEM('o031242, 16'o000000);
`MEM('o031244, 16'o000000);
`MEM('o031246, 16'o000000);
`MEM('o031250, 16'o000000);
`MEM('o031252, 16'o000000);
`MEM('o031254, 16'o000000);
`MEM('o031256, 16'o000000);
`MEM('o031260, 16'o000000);
`MEM('o031262, 16'o000000);
`MEM('o031264, 16'o000000);
`MEM('o031266, 16'o000000);
`MEM('o031270, 16'o000000);
`MEM('o031272, 16'o000000);
`MEM('o031274, 16'o000000);
`MEM('o031276, 16'o000000);
`MEM('o031300, 16'o000000);
`MEM('o031302, 16'o000000);
`MEM('o031304, 16'o000000);
`MEM('o031306, 16'o000000);
`MEM('o031310, 16'o000000);
`MEM('o031312, 16'o000000);
`MEM('o031314, 16'o000000);
`MEM('o031316, 16'o000000);
`MEM('o031320, 16'o000000);
`MEM('o031322, 16'o000000);
`MEM('o031324, 16'o000000);
`MEM('o031326, 16'o000000);
`MEM('o031330, 16'o000000);
`MEM('o031332, 16'o000000);
`MEM('o031334, 16'o000000);
`MEM('o031336, 16'o000000);
`MEM('o031340, 16'o000000);
`MEM('o031342, 16'o000000);
`MEM('o031344, 16'o000000);
`MEM('o031346, 16'o000000);
`MEM('o031350, 16'o000000);
`MEM('o031352, 16'o000000);
`MEM('o031354, 16'o000000);
`MEM('o031356, 16'o000000);
`MEM('o031360, 16'o000000);
`MEM('o031362, 16'o000000);
`MEM('o031364, 16'o000000);
`MEM('o031366, 16'o000000);
`MEM('o031370, 16'o000000);
`MEM('o031372, 16'o000000);
`MEM('o031374, 16'o000000);
`MEM('o031376, 16'o000000);
`MEM('o031400, 16'o000000);
`MEM('o031402, 16'o000000);
`MEM('o031404, 16'o000000);
`MEM('o031406, 16'o000000);
`MEM('o031410, 16'o000000);
`MEM('o031412, 16'o000000);
`MEM('o031414, 16'o000000);
`MEM('o031416, 16'o000000);
`MEM('o031420, 16'o000000);
`MEM('o031422, 16'o000000);
`MEM('o031424, 16'o000000);
`MEM('o031426, 16'o000000);
`MEM('o031430, 16'o000000);
`MEM('o031432, 16'o000000);
`MEM('o031434, 16'o000000);
`MEM('o031436, 16'o000000);
`MEM('o031440, 16'o000000);
`MEM('o031442, 16'o000000);
`MEM('o031444, 16'o000000);
`MEM('o031446, 16'o000000);
`MEM('o031450, 16'o000000);
`MEM('o031452, 16'o000000);
`MEM('o031454, 16'o000000);
`MEM('o031456, 16'o000000);
`MEM('o031460, 16'o000000);
`MEM('o031462, 16'o000000);
`MEM('o031464, 16'o000000);
`MEM('o031466, 16'o000000);
`MEM('o031470, 16'o000000);
`MEM('o031472, 16'o000000);
`MEM('o031474, 16'o000000);
`MEM('o031476, 16'o000000);
`MEM('o031500, 16'o000000);
`MEM('o031502, 16'o000000);
`MEM('o031504, 16'o000000);
`MEM('o031506, 16'o000000);
`MEM('o031510, 16'o000000);
`MEM('o031512, 16'o000000);
`MEM('o031514, 16'o000000);
`MEM('o031516, 16'o000000);
`MEM('o031520, 16'o000000);
`MEM('o031522, 16'o000000);
`MEM('o031524, 16'o000000);
`MEM('o031526, 16'o000000);
`MEM('o031530, 16'o000000);
`MEM('o031532, 16'o000000);
`MEM('o031534, 16'o000000);
`MEM('o031536, 16'o000000);
`MEM('o031540, 16'o000000);
`MEM('o031542, 16'o000000);
`MEM('o031544, 16'o000000);
`MEM('o031546, 16'o000000);
`MEM('o031550, 16'o000000);
`MEM('o031552, 16'o000000);
`MEM('o031554, 16'o000000);
`MEM('o031556, 16'o000000);
`MEM('o031560, 16'o000000);
`MEM('o031562, 16'o000000);
`MEM('o031564, 16'o000000);
`MEM('o031566, 16'o000000);
`MEM('o031570, 16'o000000);
`MEM('o031572, 16'o000000);
`MEM('o031574, 16'o000000);
`MEM('o031576, 16'o000000);
`MEM('o031600, 16'o000000);
`MEM('o031602, 16'o000000);
`MEM('o031604, 16'o000000);
`MEM('o031606, 16'o000000);
`MEM('o031610, 16'o000000);
`MEM('o031612, 16'o000000);
`MEM('o031614, 16'o000000);
`MEM('o031616, 16'o000000);
`MEM('o031620, 16'o000000);
`MEM('o031622, 16'o000000);
`MEM('o031624, 16'o000000);
`MEM('o031626, 16'o000000);
`MEM('o031630, 16'o000000);
`MEM('o031632, 16'o000000);
`MEM('o031634, 16'o000000);
`MEM('o031636, 16'o000000);
`MEM('o031640, 16'o000000);
`MEM('o031642, 16'o000000);
`MEM('o031644, 16'o000000);
`MEM('o031646, 16'o000000);
`MEM('o031650, 16'o000000);
`MEM('o031652, 16'o000000);
`MEM('o031654, 16'o000000);
`MEM('o031656, 16'o000000);
`MEM('o031660, 16'o000000);
`MEM('o031662, 16'o000000);
`MEM('o031664, 16'o000000);
`MEM('o031666, 16'o000000);
`MEM('o031670, 16'o000000);
`MEM('o031672, 16'o000000);
`MEM('o031674, 16'o000000);
`MEM('o031676, 16'o000000);
`MEM('o031700, 16'o000000);
`MEM('o031702, 16'o000000);
`MEM('o031704, 16'o000000);
`MEM('o031706, 16'o000000);
`MEM('o031710, 16'o000000);
`MEM('o031712, 16'o000000);
`MEM('o031714, 16'o000000);
`MEM('o031716, 16'o000000);
`MEM('o031720, 16'o000000);
`MEM('o031722, 16'o000000);
`MEM('o031724, 16'o000000);
`MEM('o031726, 16'o000000);
`MEM('o031730, 16'o000000);
`MEM('o031732, 16'o000000);
`MEM('o031734, 16'o000000);
`MEM('o031736, 16'o000000);
`MEM('o031740, 16'o000000);
`MEM('o031742, 16'o000000);
`MEM('o031744, 16'o000000);
`MEM('o031746, 16'o000000);
`MEM('o031750, 16'o000000);
`MEM('o031752, 16'o000000);
`MEM('o031754, 16'o000000);
`MEM('o031756, 16'o000000);
`MEM('o031760, 16'o000000);
`MEM('o031762, 16'o000000);
`MEM('o031764, 16'o000000);
`MEM('o031766, 16'o000000);
`MEM('o031770, 16'o000000);
`MEM('o031772, 16'o000000);
`MEM('o031774, 16'o000000);
`MEM('o031776, 16'o000000);
`MEM('o032000, 16'o000000);
`MEM('o032002, 16'o000000);
`MEM('o032004, 16'o000000);
`MEM('o032006, 16'o000000);
`MEM('o032010, 16'o000000);
`MEM('o032012, 16'o000000);
`MEM('o032014, 16'o000000);
`MEM('o032016, 16'o000000);
`MEM('o032020, 16'o000000);
`MEM('o032022, 16'o000000);
`MEM('o032024, 16'o000000);
`MEM('o032026, 16'o000000);
`MEM('o032030, 16'o000000);
`MEM('o032032, 16'o000000);
`MEM('o032034, 16'o000000);
`MEM('o032036, 16'o000000);
`MEM('o032040, 16'o000000);
`MEM('o032042, 16'o000000);
`MEM('o032044, 16'o000000);
`MEM('o032046, 16'o000000);
`MEM('o032050, 16'o000000);
`MEM('o032052, 16'o000000);
`MEM('o032054, 16'o000000);
`MEM('o032056, 16'o000000);
`MEM('o032060, 16'o000000);
`MEM('o032062, 16'o000000);
`MEM('o032064, 16'o000000);
`MEM('o032066, 16'o000000);
`MEM('o032070, 16'o000000);
`MEM('o032072, 16'o000000);
`MEM('o032074, 16'o000000);
`MEM('o032076, 16'o000000);
`MEM('o032100, 16'o000000);
`MEM('o032102, 16'o000000);
`MEM('o032104, 16'o000000);
`MEM('o032106, 16'o000000);
`MEM('o032110, 16'o000000);
`MEM('o032112, 16'o000000);
`MEM('o032114, 16'o000000);
`MEM('o032116, 16'o000000);
`MEM('o032120, 16'o000000);
`MEM('o032122, 16'o000000);
`MEM('o032124, 16'o000000);
`MEM('o032126, 16'o000000);
`MEM('o032130, 16'o000000);
`MEM('o032132, 16'o000000);
`MEM('o032134, 16'o000000);
`MEM('o032136, 16'o000000);
`MEM('o032140, 16'o000000);
`MEM('o032142, 16'o000000);
`MEM('o032144, 16'o000000);
`MEM('o032146, 16'o000000);
`MEM('o032150, 16'o000000);
`MEM('o032152, 16'o000000);
`MEM('o032154, 16'o000000);
`MEM('o032156, 16'o000000);
`MEM('o032160, 16'o000000);
`MEM('o032162, 16'o000000);
`MEM('o032164, 16'o000000);
`MEM('o032166, 16'o000000);
`MEM('o032170, 16'o000000);
`MEM('o032172, 16'o000000);
`MEM('o032174, 16'o000000);
`MEM('o032176, 16'o000000);
`MEM('o032200, 16'o000000);
`MEM('o032202, 16'o000000);
`MEM('o032204, 16'o000000);
`MEM('o032206, 16'o000000);
`MEM('o032210, 16'o000000);
`MEM('o032212, 16'o000000);
`MEM('o032214, 16'o000000);
`MEM('o032216, 16'o000000);
`MEM('o032220, 16'o000000);
`MEM('o032222, 16'o000000);
`MEM('o032224, 16'o000000);
`MEM('o032226, 16'o000000);
`MEM('o032230, 16'o000000);
`MEM('o032232, 16'o000000);
`MEM('o032234, 16'o000000);
`MEM('o032236, 16'o000000);
`MEM('o032240, 16'o000000);
`MEM('o032242, 16'o000000);
`MEM('o032244, 16'o000000);
`MEM('o032246, 16'o000000);
`MEM('o032250, 16'o000000);
`MEM('o032252, 16'o000000);
`MEM('o032254, 16'o000000);
`MEM('o032256, 16'o000000);
`MEM('o032260, 16'o000000);
`MEM('o032262, 16'o000000);
`MEM('o032264, 16'o000000);
`MEM('o032266, 16'o000000);
`MEM('o032270, 16'o000000);
`MEM('o032272, 16'o000000);
`MEM('o032274, 16'o000000);
`MEM('o032276, 16'o000000);
`MEM('o032300, 16'o000000);
`MEM('o032302, 16'o000000);
`MEM('o032304, 16'o000000);
`MEM('o032306, 16'o000000);
`MEM('o032310, 16'o000000);
`MEM('o032312, 16'o000000);
`MEM('o032314, 16'o000000);
`MEM('o032316, 16'o000000);
`MEM('o032320, 16'o000000);
`MEM('o032322, 16'o000000);
`MEM('o032324, 16'o000000);
`MEM('o032326, 16'o000000);
`MEM('o032330, 16'o000000);
`MEM('o032332, 16'o000000);
`MEM('o032334, 16'o000000);
`MEM('o032336, 16'o000000);
`MEM('o032340, 16'o000000);
`MEM('o032342, 16'o000000);
`MEM('o032344, 16'o000000);
`MEM('o032346, 16'o000000);
`MEM('o032350, 16'o000000);
`MEM('o032352, 16'o000000);
`MEM('o032354, 16'o000000);
`MEM('o032356, 16'o000000);
`MEM('o032360, 16'o000000);
`MEM('o032362, 16'o000000);
`MEM('o032364, 16'o000000);
`MEM('o032366, 16'o000000);
`MEM('o032370, 16'o000000);
`MEM('o032372, 16'o000000);
`MEM('o032374, 16'o000000);
`MEM('o032376, 16'o000000);
`MEM('o032400, 16'o000000);
`MEM('o032402, 16'o000000);
`MEM('o032404, 16'o000000);
`MEM('o032406, 16'o000000);
`MEM('o032410, 16'o000000);
`MEM('o032412, 16'o000000);
`MEM('o032414, 16'o000000);
`MEM('o032416, 16'o000000);
`MEM('o032420, 16'o000000);
`MEM('o032422, 16'o000000);
`MEM('o032424, 16'o000000);
`MEM('o032426, 16'o000000);
`MEM('o032430, 16'o000000);
`MEM('o032432, 16'o000000);
`MEM('o032434, 16'o000000);
`MEM('o032436, 16'o000000);
`MEM('o032440, 16'o000000);
`MEM('o032442, 16'o000000);
`MEM('o032444, 16'o000000);
`MEM('o032446, 16'o000000);
`MEM('o032450, 16'o000000);
`MEM('o032452, 16'o000000);
`MEM('o032454, 16'o000000);
`MEM('o032456, 16'o000000);
`MEM('o032460, 16'o000000);
`MEM('o032462, 16'o000000);
`MEM('o032464, 16'o000000);
`MEM('o032466, 16'o000000);
`MEM('o032470, 16'o000000);
`MEM('o032472, 16'o000000);
`MEM('o032474, 16'o000000);
`MEM('o032476, 16'o000000);
`MEM('o032500, 16'o000000);
`MEM('o032502, 16'o000000);
`MEM('o032504, 16'o000000);
`MEM('o032506, 16'o000000);
`MEM('o032510, 16'o000000);
`MEM('o032512, 16'o000000);
`MEM('o032514, 16'o000000);
`MEM('o032516, 16'o000000);
`MEM('o032520, 16'o000000);
`MEM('o032522, 16'o000000);
`MEM('o032524, 16'o000000);
`MEM('o032526, 16'o000000);
`MEM('o032530, 16'o000000);
`MEM('o032532, 16'o000000);
`MEM('o032534, 16'o000000);
`MEM('o032536, 16'o000000);
`MEM('o032540, 16'o000000);
`MEM('o032542, 16'o000000);
`MEM('o032544, 16'o000000);
`MEM('o032546, 16'o000000);
`MEM('o032550, 16'o000000);
`MEM('o032552, 16'o000000);
`MEM('o032554, 16'o000000);
`MEM('o032556, 16'o000000);
`MEM('o032560, 16'o000000);
`MEM('o032562, 16'o000000);
`MEM('o032564, 16'o000000);
`MEM('o032566, 16'o000000);
`MEM('o032570, 16'o000000);
`MEM('o032572, 16'o000000);
`MEM('o032574, 16'o000000);
`MEM('o032576, 16'o000000);
`MEM('o032600, 16'o000000);
`MEM('o032602, 16'o000000);
`MEM('o032604, 16'o000000);
`MEM('o032606, 16'o000000);
`MEM('o032610, 16'o000000);
`MEM('o032612, 16'o000000);
`MEM('o032614, 16'o000000);
`MEM('o032616, 16'o000000);
`MEM('o032620, 16'o000000);
`MEM('o032622, 16'o000000);
`MEM('o032624, 16'o000000);
`MEM('o032626, 16'o000000);
`MEM('o032630, 16'o000000);
`MEM('o032632, 16'o000000);
`MEM('o032634, 16'o000000);
`MEM('o032636, 16'o000000);
`MEM('o032640, 16'o000000);
`MEM('o032642, 16'o000000);
`MEM('o032644, 16'o000000);
`MEM('o032646, 16'o000000);
`MEM('o032650, 16'o000000);
`MEM('o032652, 16'o000000);
`MEM('o032654, 16'o000000);
`MEM('o032656, 16'o000000);
`MEM('o032660, 16'o000000);
`MEM('o032662, 16'o000000);
`MEM('o032664, 16'o000000);
`MEM('o032666, 16'o000000);
`MEM('o032670, 16'o000000);
`MEM('o032672, 16'o000000);
`MEM('o032674, 16'o000000);
`MEM('o032676, 16'o000000);
`MEM('o032700, 16'o000000);
`MEM('o032702, 16'o000000);
`MEM('o032704, 16'o000000);
`MEM('o032706, 16'o000000);
`MEM('o032710, 16'o000000);
`MEM('o032712, 16'o000000);
`MEM('o032714, 16'o000000);
`MEM('o032716, 16'o000000);
`MEM('o032720, 16'o000000);
`MEM('o032722, 16'o000000);
`MEM('o032724, 16'o000000);
`MEM('o032726, 16'o000000);
`MEM('o032730, 16'o000000);
`MEM('o032732, 16'o000000);
`MEM('o032734, 16'o000000);
`MEM('o032736, 16'o000000);
`MEM('o032740, 16'o000000);
`MEM('o032742, 16'o000000);
`MEM('o032744, 16'o000000);
`MEM('o032746, 16'o000000);
`MEM('o032750, 16'o000000);
`MEM('o032752, 16'o000000);
`MEM('o032754, 16'o000000);
`MEM('o032756, 16'o000000);
`MEM('o032760, 16'o000000);
`MEM('o032762, 16'o000000);
`MEM('o032764, 16'o000000);
`MEM('o032766, 16'o000000);
`MEM('o032770, 16'o000000);
`MEM('o032772, 16'o000000);
`MEM('o032774, 16'o000000);
`MEM('o032776, 16'o000000);
`MEM('o033000, 16'o000000);
`MEM('o033002, 16'o000000);
`MEM('o033004, 16'o000000);
`MEM('o033006, 16'o000000);
`MEM('o033010, 16'o000000);
`MEM('o033012, 16'o000000);
`MEM('o033014, 16'o000000);
`MEM('o033016, 16'o000000);
`MEM('o033020, 16'o000000);
`MEM('o033022, 16'o000000);
`MEM('o033024, 16'o000000);
`MEM('o033026, 16'o000000);
`MEM('o033030, 16'o000000);
`MEM('o033032, 16'o000000);
`MEM('o033034, 16'o000000);
`MEM('o033036, 16'o000000);
`MEM('o033040, 16'o000000);
`MEM('o033042, 16'o000000);
`MEM('o033044, 16'o000000);
`MEM('o033046, 16'o000000);
`MEM('o033050, 16'o000000);
`MEM('o033052, 16'o000000);
`MEM('o033054, 16'o000000);
`MEM('o033056, 16'o000000);
`MEM('o033060, 16'o000000);
`MEM('o033062, 16'o000000);
`MEM('o033064, 16'o000000);
`MEM('o033066, 16'o000000);
`MEM('o033070, 16'o000000);
`MEM('o033072, 16'o000000);
`MEM('o033074, 16'o000000);
`MEM('o033076, 16'o000000);
`MEM('o033100, 16'o000000);
`MEM('o033102, 16'o000000);
`MEM('o033104, 16'o000000);
`MEM('o033106, 16'o000000);
`MEM('o033110, 16'o000000);
`MEM('o033112, 16'o000000);
`MEM('o033114, 16'o000000);
`MEM('o033116, 16'o000000);
`MEM('o033120, 16'o000000);
`MEM('o033122, 16'o000000);
`MEM('o033124, 16'o000000);
`MEM('o033126, 16'o000000);
`MEM('o033130, 16'o000000);
`MEM('o033132, 16'o000000);
`MEM('o033134, 16'o000000);
`MEM('o033136, 16'o000000);
`MEM('o033140, 16'o000000);
`MEM('o033142, 16'o000000);
`MEM('o033144, 16'o000000);
`MEM('o033146, 16'o000000);
`MEM('o033150, 16'o000000);
`MEM('o033152, 16'o000000);
`MEM('o033154, 16'o000000);
`MEM('o033156, 16'o000000);
`MEM('o033160, 16'o000000);
`MEM('o033162, 16'o000000);
`MEM('o033164, 16'o000000);
`MEM('o033166, 16'o000000);
`MEM('o033170, 16'o000000);
`MEM('o033172, 16'o000000);
`MEM('o033174, 16'o000000);
`MEM('o033176, 16'o000000);
`MEM('o033200, 16'o000000);
`MEM('o033202, 16'o000000);
`MEM('o033204, 16'o000000);
`MEM('o033206, 16'o000000);
`MEM('o033210, 16'o000000);
`MEM('o033212, 16'o000000);
`MEM('o033214, 16'o000000);
`MEM('o033216, 16'o000000);
`MEM('o033220, 16'o000000);
`MEM('o033222, 16'o000000);
`MEM('o033224, 16'o000000);
`MEM('o033226, 16'o000000);
`MEM('o033230, 16'o000000);
`MEM('o033232, 16'o000000);
`MEM('o033234, 16'o000000);
`MEM('o033236, 16'o000000);
`MEM('o033240, 16'o000000);
`MEM('o033242, 16'o000000);
`MEM('o033244, 16'o000000);
`MEM('o033246, 16'o000000);
`MEM('o033250, 16'o000000);
`MEM('o033252, 16'o000000);
`MEM('o033254, 16'o000000);
`MEM('o033256, 16'o000000);
`MEM('o033260, 16'o000000);
`MEM('o033262, 16'o000000);
`MEM('o033264, 16'o000000);
`MEM('o033266, 16'o000000);
`MEM('o033270, 16'o000000);
`MEM('o033272, 16'o000000);
`MEM('o033274, 16'o000000);
`MEM('o033276, 16'o000000);
`MEM('o033300, 16'o000000);
`MEM('o033302, 16'o000000);
`MEM('o033304, 16'o000000);
`MEM('o033306, 16'o000000);
`MEM('o033310, 16'o000000);
`MEM('o033312, 16'o000000);
`MEM('o033314, 16'o000000);
`MEM('o033316, 16'o000000);
`MEM('o033320, 16'o000000);
`MEM('o033322, 16'o000000);
`MEM('o033324, 16'o000000);
`MEM('o033326, 16'o000000);
`MEM('o033330, 16'o000000);
`MEM('o033332, 16'o000000);
`MEM('o033334, 16'o000000);
`MEM('o033336, 16'o000000);
`MEM('o033340, 16'o000000);
`MEM('o033342, 16'o000000);
`MEM('o033344, 16'o000000);
`MEM('o033346, 16'o000000);
`MEM('o033350, 16'o000000);
`MEM('o033352, 16'o000000);
`MEM('o033354, 16'o000000);
`MEM('o033356, 16'o000000);
`MEM('o033360, 16'o000000);
`MEM('o033362, 16'o000000);
`MEM('o033364, 16'o000000);
`MEM('o033366, 16'o000000);
`MEM('o033370, 16'o000000);
`MEM('o033372, 16'o000000);
`MEM('o033374, 16'o000000);
`MEM('o033376, 16'o000000);
`MEM('o033400, 16'o000000);
`MEM('o033402, 16'o000000);
`MEM('o033404, 16'o000000);
`MEM('o033406, 16'o000000);
`MEM('o033410, 16'o000000);
`MEM('o033412, 16'o000000);
`MEM('o033414, 16'o000000);
`MEM('o033416, 16'o000000);
`MEM('o033420, 16'o000000);
`MEM('o033422, 16'o000000);
`MEM('o033424, 16'o000000);
`MEM('o033426, 16'o000000);
`MEM('o033430, 16'o000000);
`MEM('o033432, 16'o000000);
`MEM('o033434, 16'o000000);
`MEM('o033436, 16'o000000);
`MEM('o033440, 16'o000000);
`MEM('o033442, 16'o000000);
`MEM('o033444, 16'o000000);
`MEM('o033446, 16'o000000);
`MEM('o033450, 16'o000000);
`MEM('o033452, 16'o000000);
`MEM('o033454, 16'o000000);
`MEM('o033456, 16'o000000);
`MEM('o033460, 16'o000000);
`MEM('o033462, 16'o000000);
`MEM('o033464, 16'o000000);
`MEM('o033466, 16'o000000);
`MEM('o033470, 16'o000000);
`MEM('o033472, 16'o000000);
`MEM('o033474, 16'o000000);
`MEM('o033476, 16'o000000);
`MEM('o033500, 16'o000000);
`MEM('o033502, 16'o000000);
`MEM('o033504, 16'o000000);
`MEM('o033506, 16'o000000);
`MEM('o033510, 16'o000000);
`MEM('o033512, 16'o000000);
`MEM('o033514, 16'o000000);
`MEM('o033516, 16'o000000);
`MEM('o033520, 16'o000000);
`MEM('o033522, 16'o000000);
`MEM('o033524, 16'o000000);
`MEM('o033526, 16'o000000);
`MEM('o033530, 16'o000000);
`MEM('o033532, 16'o000000);
`MEM('o033534, 16'o000000);
`MEM('o033536, 16'o000000);
`MEM('o033540, 16'o000000);
`MEM('o033542, 16'o000000);
`MEM('o033544, 16'o000000);
`MEM('o033546, 16'o000000);
`MEM('o033550, 16'o000000);
`MEM('o033552, 16'o000000);
`MEM('o033554, 16'o000000);
`MEM('o033556, 16'o000000);
`MEM('o033560, 16'o000000);
`MEM('o033562, 16'o000000);
`MEM('o033564, 16'o000000);
`MEM('o033566, 16'o000000);
`MEM('o033570, 16'o000000);
`MEM('o033572, 16'o000000);
`MEM('o033574, 16'o000000);
`MEM('o033576, 16'o000000);
`MEM('o033600, 16'o000000);
`MEM('o033602, 16'o000000);
`MEM('o033604, 16'o000000);
`MEM('o033606, 16'o000000);
`MEM('o033610, 16'o000000);
`MEM('o033612, 16'o000000);
`MEM('o033614, 16'o000000);
`MEM('o033616, 16'o000000);
`MEM('o033620, 16'o000000);
`MEM('o033622, 16'o000000);
`MEM('o033624, 16'o000000);
`MEM('o033626, 16'o000000);
`MEM('o033630, 16'o000000);
`MEM('o033632, 16'o000000);
`MEM('o033634, 16'o000000);
`MEM('o033636, 16'o000000);
`MEM('o033640, 16'o000000);
`MEM('o033642, 16'o000000);
`MEM('o033644, 16'o000000);
`MEM('o033646, 16'o000000);
`MEM('o033650, 16'o000000);
`MEM('o033652, 16'o000000);
`MEM('o033654, 16'o000000);
`MEM('o033656, 16'o000000);
`MEM('o033660, 16'o000000);
`MEM('o033662, 16'o000000);
`MEM('o033664, 16'o000000);
`MEM('o033666, 16'o000000);
`MEM('o033670, 16'o000000);
`MEM('o033672, 16'o000000);
`MEM('o033674, 16'o000000);
`MEM('o033676, 16'o000000);
`MEM('o033700, 16'o000000);
`MEM('o033702, 16'o000000);
`MEM('o033704, 16'o000000);
`MEM('o033706, 16'o000000);
`MEM('o033710, 16'o000000);
`MEM('o033712, 16'o000000);
`MEM('o033714, 16'o000000);
`MEM('o033716, 16'o000000);
`MEM('o033720, 16'o000000);
`MEM('o033722, 16'o000000);
`MEM('o033724, 16'o000000);
`MEM('o033726, 16'o000000);
`MEM('o033730, 16'o000000);
`MEM('o033732, 16'o000000);
`MEM('o033734, 16'o000000);
`MEM('o033736, 16'o000000);
`MEM('o033740, 16'o000000);
`MEM('o033742, 16'o000000);
`MEM('o033744, 16'o000000);
`MEM('o033746, 16'o000000);
`MEM('o033750, 16'o000000);
`MEM('o033752, 16'o000000);
`MEM('o033754, 16'o000000);
`MEM('o033756, 16'o000000);
`MEM('o033760, 16'o000000);
`MEM('o033762, 16'o000000);
`MEM('o033764, 16'o000000);
`MEM('o033766, 16'o000000);
`MEM('o033770, 16'o000000);
`MEM('o033772, 16'o000000);
`MEM('o033774, 16'o000000);
`MEM('o033776, 16'o000000);
`MEM('o034000, 16'o000000);
`MEM('o034002, 16'o000000);
`MEM('o034004, 16'o000000);
`MEM('o034006, 16'o000000);
`MEM('o034010, 16'o000000);
`MEM('o034012, 16'o000000);
`MEM('o034014, 16'o000000);
`MEM('o034016, 16'o000000);
`MEM('o034020, 16'o000000);
`MEM('o034022, 16'o000000);
`MEM('o034024, 16'o000000);
`MEM('o034026, 16'o000000);
`MEM('o034030, 16'o000000);
`MEM('o034032, 16'o000000);
`MEM('o034034, 16'o000000);
`MEM('o034036, 16'o000000);
`MEM('o034040, 16'o000000);
`MEM('o034042, 16'o000000);
`MEM('o034044, 16'o000000);
`MEM('o034046, 16'o000000);
`MEM('o034050, 16'o000000);
`MEM('o034052, 16'o000000);
`MEM('o034054, 16'o000000);
`MEM('o034056, 16'o000000);
`MEM('o034060, 16'o000000);
`MEM('o034062, 16'o000000);
`MEM('o034064, 16'o000000);
`MEM('o034066, 16'o000000);
`MEM('o034070, 16'o000000);
`MEM('o034072, 16'o000000);
`MEM('o034074, 16'o000000);
`MEM('o034076, 16'o000000);
`MEM('o034100, 16'o000000);
`MEM('o034102, 16'o000000);
`MEM('o034104, 16'o000000);
`MEM('o034106, 16'o000000);
`MEM('o034110, 16'o000000);
`MEM('o034112, 16'o000000);
`MEM('o034114, 16'o000000);
`MEM('o034116, 16'o000000);
`MEM('o034120, 16'o000000);
`MEM('o034122, 16'o000000);
`MEM('o034124, 16'o000000);
`MEM('o034126, 16'o000000);
`MEM('o034130, 16'o000000);
`MEM('o034132, 16'o000000);
`MEM('o034134, 16'o000000);
`MEM('o034136, 16'o000000);
`MEM('o034140, 16'o000000);
`MEM('o034142, 16'o000000);
`MEM('o034144, 16'o000000);
`MEM('o034146, 16'o000000);
`MEM('o034150, 16'o000000);
`MEM('o034152, 16'o000000);
`MEM('o034154, 16'o000000);
`MEM('o034156, 16'o000000);
`MEM('o034160, 16'o000000);
`MEM('o034162, 16'o000000);
`MEM('o034164, 16'o000000);
`MEM('o034166, 16'o000000);
`MEM('o034170, 16'o000000);
`MEM('o034172, 16'o000000);
`MEM('o034174, 16'o000000);
`MEM('o034176, 16'o000000);
`MEM('o034200, 16'o000000);
`MEM('o034202, 16'o000000);
`MEM('o034204, 16'o000000);
`MEM('o034206, 16'o000000);
`MEM('o034210, 16'o000000);
`MEM('o034212, 16'o000000);
`MEM('o034214, 16'o000000);
`MEM('o034216, 16'o000000);
`MEM('o034220, 16'o000000);
`MEM('o034222, 16'o000000);
`MEM('o034224, 16'o000000);
`MEM('o034226, 16'o000000);
`MEM('o034230, 16'o000000);
`MEM('o034232, 16'o000000);
`MEM('o034234, 16'o000000);
`MEM('o034236, 16'o000000);
`MEM('o034240, 16'o000000);
`MEM('o034242, 16'o000000);
`MEM('o034244, 16'o000000);
`MEM('o034246, 16'o000000);
`MEM('o034250, 16'o000000);
`MEM('o034252, 16'o000000);
`MEM('o034254, 16'o000000);
`MEM('o034256, 16'o000000);
`MEM('o034260, 16'o000000);
`MEM('o034262, 16'o000000);
`MEM('o034264, 16'o000000);
`MEM('o034266, 16'o000000);
`MEM('o034270, 16'o000000);
`MEM('o034272, 16'o000000);
`MEM('o034274, 16'o000000);
`MEM('o034276, 16'o000000);
`MEM('o034300, 16'o000000);
`MEM('o034302, 16'o000000);
`MEM('o034304, 16'o000000);
`MEM('o034306, 16'o000000);
`MEM('o034310, 16'o000000);
`MEM('o034312, 16'o000000);
`MEM('o034314, 16'o000000);
`MEM('o034316, 16'o000000);
`MEM('o034320, 16'o000000);
`MEM('o034322, 16'o000000);
`MEM('o034324, 16'o000000);
`MEM('o034326, 16'o000000);
`MEM('o034330, 16'o000000);
`MEM('o034332, 16'o000000);
`MEM('o034334, 16'o000000);
`MEM('o034336, 16'o000000);
`MEM('o034340, 16'o000000);
`MEM('o034342, 16'o000000);
`MEM('o034344, 16'o000000);
`MEM('o034346, 16'o000000);
`MEM('o034350, 16'o000000);
`MEM('o034352, 16'o000000);
`MEM('o034354, 16'o000000);
`MEM('o034356, 16'o000000);
`MEM('o034360, 16'o000000);
`MEM('o034362, 16'o000000);
`MEM('o034364, 16'o000000);
`MEM('o034366, 16'o000000);
`MEM('o034370, 16'o000000);
`MEM('o034372, 16'o000000);
`MEM('o034374, 16'o000000);
`MEM('o034376, 16'o000000);
`MEM('o034400, 16'o000000);
`MEM('o034402, 16'o000000);
`MEM('o034404, 16'o000000);
`MEM('o034406, 16'o000000);
`MEM('o034410, 16'o000000);
`MEM('o034412, 16'o000000);
`MEM('o034414, 16'o000000);
`MEM('o034416, 16'o000000);
`MEM('o034420, 16'o000000);
`MEM('o034422, 16'o000000);
`MEM('o034424, 16'o000000);
`MEM('o034426, 16'o000000);
`MEM('o034430, 16'o000000);
`MEM('o034432, 16'o000000);
`MEM('o034434, 16'o000000);
`MEM('o034436, 16'o000000);
`MEM('o034440, 16'o000000);
`MEM('o034442, 16'o000000);
`MEM('o034444, 16'o000000);
`MEM('o034446, 16'o000000);
`MEM('o034450, 16'o000000);
`MEM('o034452, 16'o000000);
`MEM('o034454, 16'o000000);
`MEM('o034456, 16'o000000);
`MEM('o034460, 16'o000000);
`MEM('o034462, 16'o000000);
`MEM('o034464, 16'o000000);
`MEM('o034466, 16'o000000);
`MEM('o034470, 16'o000000);
`MEM('o034472, 16'o000000);
`MEM('o034474, 16'o000000);
`MEM('o034476, 16'o000000);
`MEM('o034500, 16'o000000);
`MEM('o034502, 16'o000000);
`MEM('o034504, 16'o000000);
`MEM('o034506, 16'o000000);
`MEM('o034510, 16'o000000);
`MEM('o034512, 16'o000000);
`MEM('o034514, 16'o000000);
`MEM('o034516, 16'o000000);
`MEM('o034520, 16'o000000);
`MEM('o034522, 16'o000000);
`MEM('o034524, 16'o000000);
`MEM('o034526, 16'o000000);
`MEM('o034530, 16'o000000);
`MEM('o034532, 16'o000000);
`MEM('o034534, 16'o000000);
`MEM('o034536, 16'o000000);
`MEM('o034540, 16'o000000);
`MEM('o034542, 16'o000000);
`MEM('o034544, 16'o000000);
`MEM('o034546, 16'o000000);
`MEM('o034550, 16'o000000);
`MEM('o034552, 16'o000000);
`MEM('o034554, 16'o000000);
`MEM('o034556, 16'o000000);
`MEM('o034560, 16'o000000);
`MEM('o034562, 16'o000000);
`MEM('o034564, 16'o000000);
`MEM('o034566, 16'o000000);
`MEM('o034570, 16'o000000);
`MEM('o034572, 16'o000000);
`MEM('o034574, 16'o000000);
`MEM('o034576, 16'o000000);
`MEM('o034600, 16'o000000);
`MEM('o034602, 16'o000000);
`MEM('o034604, 16'o000000);
`MEM('o034606, 16'o000000);
`MEM('o034610, 16'o000000);
`MEM('o034612, 16'o000000);
`MEM('o034614, 16'o000000);
`MEM('o034616, 16'o000000);
`MEM('o034620, 16'o000000);
`MEM('o034622, 16'o000000);
`MEM('o034624, 16'o000000);
`MEM('o034626, 16'o000000);
`MEM('o034630, 16'o000000);
`MEM('o034632, 16'o000000);
`MEM('o034634, 16'o000000);
`MEM('o034636, 16'o000000);
`MEM('o034640, 16'o000000);
`MEM('o034642, 16'o000000);
`MEM('o034644, 16'o000000);
`MEM('o034646, 16'o000000);
`MEM('o034650, 16'o000000);
`MEM('o034652, 16'o000000);
`MEM('o034654, 16'o000000);
`MEM('o034656, 16'o000000);
`MEM('o034660, 16'o000000);
`MEM('o034662, 16'o000000);
`MEM('o034664, 16'o000000);
`MEM('o034666, 16'o000000);
`MEM('o034670, 16'o000000);
`MEM('o034672, 16'o000000);
`MEM('o034674, 16'o000000);
`MEM('o034676, 16'o000000);
`MEM('o034700, 16'o000000);
`MEM('o034702, 16'o000000);
`MEM('o034704, 16'o000000);
`MEM('o034706, 16'o000000);
`MEM('o034710, 16'o000000);
`MEM('o034712, 16'o000000);
`MEM('o034714, 16'o000000);
`MEM('o034716, 16'o000000);
`MEM('o034720, 16'o000000);
`MEM('o034722, 16'o000000);
`MEM('o034724, 16'o000000);
`MEM('o034726, 16'o000000);
`MEM('o034730, 16'o000000);
`MEM('o034732, 16'o000000);
`MEM('o034734, 16'o000000);
`MEM('o034736, 16'o000000);
`MEM('o034740, 16'o000000);
`MEM('o034742, 16'o000000);
`MEM('o034744, 16'o000000);
`MEM('o034746, 16'o000000);
`MEM('o034750, 16'o000000);
`MEM('o034752, 16'o000000);
`MEM('o034754, 16'o000000);
`MEM('o034756, 16'o000000);
`MEM('o034760, 16'o000000);
`MEM('o034762, 16'o000000);
`MEM('o034764, 16'o000000);
`MEM('o034766, 16'o000000);
`MEM('o034770, 16'o000000);
`MEM('o034772, 16'o000000);
`MEM('o034774, 16'o000000);
`MEM('o034776, 16'o000000);
`MEM('o035000, 16'o000000);
`MEM('o035002, 16'o000000);
`MEM('o035004, 16'o000000);
`MEM('o035006, 16'o000000);
`MEM('o035010, 16'o000000);
`MEM('o035012, 16'o000000);
`MEM('o035014, 16'o000000);
`MEM('o035016, 16'o000000);
`MEM('o035020, 16'o000000);
`MEM('o035022, 16'o000000);
`MEM('o035024, 16'o000000);
`MEM('o035026, 16'o000000);
`MEM('o035030, 16'o000000);
`MEM('o035032, 16'o000000);
`MEM('o035034, 16'o000000);
`MEM('o035036, 16'o000000);
`MEM('o035040, 16'o000000);
`MEM('o035042, 16'o000000);
`MEM('o035044, 16'o000000);
`MEM('o035046, 16'o000000);
`MEM('o035050, 16'o000000);
`MEM('o035052, 16'o000000);
`MEM('o035054, 16'o000000);
`MEM('o035056, 16'o000000);
`MEM('o035060, 16'o000000);
`MEM('o035062, 16'o000000);
`MEM('o035064, 16'o000000);
`MEM('o035066, 16'o000000);
`MEM('o035070, 16'o000000);
`MEM('o035072, 16'o000000);
`MEM('o035074, 16'o000000);
`MEM('o035076, 16'o000000);
`MEM('o035100, 16'o000000);
`MEM('o035102, 16'o000000);
`MEM('o035104, 16'o000000);
`MEM('o035106, 16'o000000);
`MEM('o035110, 16'o000000);
`MEM('o035112, 16'o000000);
`MEM('o035114, 16'o000000);
`MEM('o035116, 16'o000000);
`MEM('o035120, 16'o000000);
`MEM('o035122, 16'o000000);
`MEM('o035124, 16'o000000);
`MEM('o035126, 16'o000000);
`MEM('o035130, 16'o000000);
`MEM('o035132, 16'o000000);
`MEM('o035134, 16'o000000);
`MEM('o035136, 16'o000000);
`MEM('o035140, 16'o000000);
`MEM('o035142, 16'o000000);
`MEM('o035144, 16'o000000);
`MEM('o035146, 16'o000000);
`MEM('o035150, 16'o000000);
`MEM('o035152, 16'o000000);
`MEM('o035154, 16'o000000);
`MEM('o035156, 16'o000000);
`MEM('o035160, 16'o000000);
`MEM('o035162, 16'o000000);
`MEM('o035164, 16'o000000);
`MEM('o035166, 16'o000000);
`MEM('o035170, 16'o000000);
`MEM('o035172, 16'o000000);
`MEM('o035174, 16'o000000);
`MEM('o035176, 16'o000000);
`MEM('o035200, 16'o000000);
`MEM('o035202, 16'o000000);
`MEM('o035204, 16'o000000);
`MEM('o035206, 16'o000000);
`MEM('o035210, 16'o000000);
`MEM('o035212, 16'o000000);
`MEM('o035214, 16'o000000);
`MEM('o035216, 16'o000000);
`MEM('o035220, 16'o000000);
`MEM('o035222, 16'o000000);
`MEM('o035224, 16'o000000);
`MEM('o035226, 16'o000000);
`MEM('o035230, 16'o000000);
`MEM('o035232, 16'o000000);
`MEM('o035234, 16'o000000);
`MEM('o035236, 16'o000000);
`MEM('o035240, 16'o000000);
`MEM('o035242, 16'o000000);
`MEM('o035244, 16'o000000);
`MEM('o035246, 16'o000000);
`MEM('o035250, 16'o000000);
`MEM('o035252, 16'o000000);
`MEM('o035254, 16'o000000);
`MEM('o035256, 16'o000000);
`MEM('o035260, 16'o000000);
`MEM('o035262, 16'o000000);
`MEM('o035264, 16'o000000);
`MEM('o035266, 16'o000000);
`MEM('o035270, 16'o000000);
`MEM('o035272, 16'o000000);
`MEM('o035274, 16'o000000);
`MEM('o035276, 16'o000000);
`MEM('o035300, 16'o000000);
`MEM('o035302, 16'o000000);
`MEM('o035304, 16'o000000);
`MEM('o035306, 16'o000000);
`MEM('o035310, 16'o000000);
`MEM('o035312, 16'o000000);
`MEM('o035314, 16'o000000);
`MEM('o035316, 16'o000000);
`MEM('o035320, 16'o000000);
`MEM('o035322, 16'o000000);
`MEM('o035324, 16'o000000);
`MEM('o035326, 16'o000000);
`MEM('o035330, 16'o000000);
`MEM('o035332, 16'o000000);
`MEM('o035334, 16'o000000);
`MEM('o035336, 16'o000000);
`MEM('o035340, 16'o000000);
`MEM('o035342, 16'o000000);
`MEM('o035344, 16'o000000);
`MEM('o035346, 16'o000000);
`MEM('o035350, 16'o000000);
`MEM('o035352, 16'o000000);
`MEM('o035354, 16'o000000);
`MEM('o035356, 16'o000000);
`MEM('o035360, 16'o000000);
`MEM('o035362, 16'o000000);
`MEM('o035364, 16'o000000);
`MEM('o035366, 16'o000000);
`MEM('o035370, 16'o000000);
`MEM('o035372, 16'o000000);
`MEM('o035374, 16'o000000);
`MEM('o035376, 16'o000000);
`MEM('o035400, 16'o000000);
`MEM('o035402, 16'o000000);
`MEM('o035404, 16'o000000);
`MEM('o035406, 16'o000000);
`MEM('o035410, 16'o000000);
`MEM('o035412, 16'o000000);
`MEM('o035414, 16'o000000);
`MEM('o035416, 16'o000000);
`MEM('o035420, 16'o000000);
`MEM('o035422, 16'o000000);
`MEM('o035424, 16'o000000);
`MEM('o035426, 16'o000000);
`MEM('o035430, 16'o000000);
`MEM('o035432, 16'o000000);
`MEM('o035434, 16'o000000);
`MEM('o035436, 16'o000000);
`MEM('o035440, 16'o000000);
`MEM('o035442, 16'o000000);
`MEM('o035444, 16'o000000);
`MEM('o035446, 16'o000000);
`MEM('o035450, 16'o000000);
`MEM('o035452, 16'o000000);
`MEM('o035454, 16'o000000);
`MEM('o035456, 16'o000000);
`MEM('o035460, 16'o000000);
`MEM('o035462, 16'o000000);
`MEM('o035464, 16'o000000);
`MEM('o035466, 16'o000000);
`MEM('o035470, 16'o000000);
`MEM('o035472, 16'o000000);
`MEM('o035474, 16'o000000);
`MEM('o035476, 16'o000000);
`MEM('o035500, 16'o000000);
`MEM('o035502, 16'o000000);
`MEM('o035504, 16'o000000);
`MEM('o035506, 16'o000000);
`MEM('o035510, 16'o000000);
`MEM('o035512, 16'o000000);
`MEM('o035514, 16'o000000);
`MEM('o035516, 16'o000000);
`MEM('o035520, 16'o000000);
`MEM('o035522, 16'o000000);
`MEM('o035524, 16'o000000);
`MEM('o035526, 16'o000000);
`MEM('o035530, 16'o000000);
`MEM('o035532, 16'o000000);
`MEM('o035534, 16'o000000);
`MEM('o035536, 16'o000000);
`MEM('o035540, 16'o000000);
`MEM('o035542, 16'o000000);
`MEM('o035544, 16'o000000);
`MEM('o035546, 16'o000000);
`MEM('o035550, 16'o000000);
`MEM('o035552, 16'o000000);
`MEM('o035554, 16'o000000);
`MEM('o035556, 16'o000000);
`MEM('o035560, 16'o000000);
`MEM('o035562, 16'o000000);
`MEM('o035564, 16'o000000);
`MEM('o035566, 16'o000000);
`MEM('o035570, 16'o000000);
`MEM('o035572, 16'o000000);
`MEM('o035574, 16'o000000);
`MEM('o035576, 16'o000000);
`MEM('o035600, 16'o000000);
`MEM('o035602, 16'o000000);
`MEM('o035604, 16'o000000);
`MEM('o035606, 16'o000000);
`MEM('o035610, 16'o000000);
`MEM('o035612, 16'o000000);
`MEM('o035614, 16'o000000);
`MEM('o035616, 16'o000000);
`MEM('o035620, 16'o000000);
`MEM('o035622, 16'o000000);
`MEM('o035624, 16'o000000);
`MEM('o035626, 16'o000000);
`MEM('o035630, 16'o000000);
`MEM('o035632, 16'o000000);
`MEM('o035634, 16'o000000);
`MEM('o035636, 16'o000000);
`MEM('o035640, 16'o000000);
`MEM('o035642, 16'o000000);
`MEM('o035644, 16'o000000);
`MEM('o035646, 16'o000000);
`MEM('o035650, 16'o000000);
`MEM('o035652, 16'o000000);
`MEM('o035654, 16'o000000);
`MEM('o035656, 16'o000000);
`MEM('o035660, 16'o000000);
`MEM('o035662, 16'o000000);
`MEM('o035664, 16'o000000);
`MEM('o035666, 16'o000000);
`MEM('o035670, 16'o000000);
`MEM('o035672, 16'o000000);
`MEM('o035674, 16'o000000);
`MEM('o035676, 16'o000000);
`MEM('o035700, 16'o000000);
`MEM('o035702, 16'o000000);
`MEM('o035704, 16'o000000);
`MEM('o035706, 16'o000000);
`MEM('o035710, 16'o000000);
`MEM('o035712, 16'o000000);
`MEM('o035714, 16'o000000);
`MEM('o035716, 16'o000000);
`MEM('o035720, 16'o000000);
`MEM('o035722, 16'o000000);
`MEM('o035724, 16'o000000);
`MEM('o035726, 16'o000000);
`MEM('o035730, 16'o000000);
`MEM('o035732, 16'o000000);
`MEM('o035734, 16'o000000);
`MEM('o035736, 16'o000000);
`MEM('o035740, 16'o000000);
`MEM('o035742, 16'o000000);
`MEM('o035744, 16'o000000);
`MEM('o035746, 16'o000000);
`MEM('o035750, 16'o000000);
`MEM('o035752, 16'o000000);
`MEM('o035754, 16'o000000);
`MEM('o035756, 16'o000000);
`MEM('o035760, 16'o000000);
`MEM('o035762, 16'o000000);
`MEM('o035764, 16'o000000);
`MEM('o035766, 16'o000000);
`MEM('o035770, 16'o000000);
`MEM('o035772, 16'o000000);
`MEM('o035774, 16'o000000);
`MEM('o035776, 16'o000000);
`MEM('o036000, 16'o000000);
`MEM('o036002, 16'o000000);
`MEM('o036004, 16'o000000);
`MEM('o036006, 16'o000000);
`MEM('o036010, 16'o000000);
`MEM('o036012, 16'o000000);
`MEM('o036014, 16'o000000);
`MEM('o036016, 16'o000000);
`MEM('o036020, 16'o000000);
`MEM('o036022, 16'o000000);
`MEM('o036024, 16'o000000);
`MEM('o036026, 16'o000000);
`MEM('o036030, 16'o000000);
`MEM('o036032, 16'o000000);
`MEM('o036034, 16'o000000);
`MEM('o036036, 16'o000000);
`MEM('o036040, 16'o000000);
`MEM('o036042, 16'o000000);
`MEM('o036044, 16'o000000);
`MEM('o036046, 16'o000000);
`MEM('o036050, 16'o000000);
`MEM('o036052, 16'o000000);
`MEM('o036054, 16'o000000);
`MEM('o036056, 16'o000000);
`MEM('o036060, 16'o000000);
`MEM('o036062, 16'o000000);
`MEM('o036064, 16'o000000);
`MEM('o036066, 16'o000000);
`MEM('o036070, 16'o000000);
`MEM('o036072, 16'o000000);
`MEM('o036074, 16'o000000);
`MEM('o036076, 16'o000000);
`MEM('o036100, 16'o000000);
`MEM('o036102, 16'o000000);
`MEM('o036104, 16'o000000);
`MEM('o036106, 16'o000000);
`MEM('o036110, 16'o000000);
`MEM('o036112, 16'o000000);
`MEM('o036114, 16'o000000);
`MEM('o036116, 16'o000000);
`MEM('o036120, 16'o000000);
`MEM('o036122, 16'o000000);
`MEM('o036124, 16'o000000);
`MEM('o036126, 16'o000000);
`MEM('o036130, 16'o000000);
`MEM('o036132, 16'o000000);
`MEM('o036134, 16'o000000);
`MEM('o036136, 16'o000000);
`MEM('o036140, 16'o000000);
`MEM('o036142, 16'o000000);
`MEM('o036144, 16'o000000);
`MEM('o036146, 16'o000000);
`MEM('o036150, 16'o000000);
`MEM('o036152, 16'o000000);
`MEM('o036154, 16'o000000);
`MEM('o036156, 16'o000000);
`MEM('o036160, 16'o000000);
`MEM('o036162, 16'o000000);
`MEM('o036164, 16'o000000);
`MEM('o036166, 16'o000000);
`MEM('o036170, 16'o000000);
`MEM('o036172, 16'o000000);
`MEM('o036174, 16'o000000);
`MEM('o036176, 16'o000000);
`MEM('o036200, 16'o000000);
`MEM('o036202, 16'o000000);
`MEM('o036204, 16'o000000);
`MEM('o036206, 16'o000000);
`MEM('o036210, 16'o000000);
`MEM('o036212, 16'o000000);
`MEM('o036214, 16'o000000);
`MEM('o036216, 16'o000000);
`MEM('o036220, 16'o000000);
`MEM('o036222, 16'o000000);
`MEM('o036224, 16'o000000);
`MEM('o036226, 16'o000000);
`MEM('o036230, 16'o000000);
`MEM('o036232, 16'o000000);
`MEM('o036234, 16'o000000);
`MEM('o036236, 16'o000000);
`MEM('o036240, 16'o000000);
`MEM('o036242, 16'o000000);
`MEM('o036244, 16'o000000);
`MEM('o036246, 16'o000000);
`MEM('o036250, 16'o000000);
`MEM('o036252, 16'o000000);
`MEM('o036254, 16'o000000);
`MEM('o036256, 16'o000000);
`MEM('o036260, 16'o000000);
`MEM('o036262, 16'o000000);
`MEM('o036264, 16'o000000);
`MEM('o036266, 16'o000000);
`MEM('o036270, 16'o000000);
`MEM('o036272, 16'o000000);
`MEM('o036274, 16'o000000);
`MEM('o036276, 16'o000000);
`MEM('o036300, 16'o000000);
`MEM('o036302, 16'o000000);
`MEM('o036304, 16'o000000);
`MEM('o036306, 16'o000000);
`MEM('o036310, 16'o000000);
`MEM('o036312, 16'o000000);
`MEM('o036314, 16'o000000);
`MEM('o036316, 16'o000000);
`MEM('o036320, 16'o000000);
`MEM('o036322, 16'o000000);
`MEM('o036324, 16'o000000);
`MEM('o036326, 16'o000000);
`MEM('o036330, 16'o000000);
`MEM('o036332, 16'o000000);
`MEM('o036334, 16'o000000);
`MEM('o036336, 16'o000000);
`MEM('o036340, 16'o000000);
`MEM('o036342, 16'o000000);
`MEM('o036344, 16'o000000);
`MEM('o036346, 16'o000000);
`MEM('o036350, 16'o000000);
`MEM('o036352, 16'o000000);
`MEM('o036354, 16'o000000);
`MEM('o036356, 16'o000000);
`MEM('o036360, 16'o000000);
`MEM('o036362, 16'o000000);
`MEM('o036364, 16'o000000);
`MEM('o036366, 16'o000000);
`MEM('o036370, 16'o000000);
`MEM('o036372, 16'o000000);
`MEM('o036374, 16'o000000);
`MEM('o036376, 16'o000000);
`MEM('o036400, 16'o000000);
`MEM('o036402, 16'o000000);
`MEM('o036404, 16'o000000);
`MEM('o036406, 16'o000000);
`MEM('o036410, 16'o000000);
`MEM('o036412, 16'o000000);
`MEM('o036414, 16'o000000);
`MEM('o036416, 16'o000000);
`MEM('o036420, 16'o000000);
`MEM('o036422, 16'o000000);
`MEM('o036424, 16'o000000);
`MEM('o036426, 16'o000000);
`MEM('o036430, 16'o000000);
`MEM('o036432, 16'o000000);
`MEM('o036434, 16'o000000);
`MEM('o036436, 16'o000000);
`MEM('o036440, 16'o000000);
`MEM('o036442, 16'o000000);
`MEM('o036444, 16'o000000);
`MEM('o036446, 16'o000000);
`MEM('o036450, 16'o000000);
`MEM('o036452, 16'o000000);
`MEM('o036454, 16'o000000);
`MEM('o036456, 16'o000000);
`MEM('o036460, 16'o000000);
`MEM('o036462, 16'o000000);
`MEM('o036464, 16'o000000);
`MEM('o036466, 16'o000000);
`MEM('o036470, 16'o000000);
`MEM('o036472, 16'o000000);
`MEM('o036474, 16'o000000);
`MEM('o036476, 16'o000000);
`MEM('o036500, 16'o000000);
`MEM('o036502, 16'o000000);
`MEM('o036504, 16'o000000);
`MEM('o036506, 16'o000000);
`MEM('o036510, 16'o000000);
`MEM('o036512, 16'o000000);
`MEM('o036514, 16'o000000);
`MEM('o036516, 16'o000000);
`MEM('o036520, 16'o000000);
`MEM('o036522, 16'o000000);
`MEM('o036524, 16'o000000);
`MEM('o036526, 16'o000000);
`MEM('o036530, 16'o000000);
`MEM('o036532, 16'o000000);
`MEM('o036534, 16'o000000);
`MEM('o036536, 16'o000000);
`MEM('o036540, 16'o000000);
`MEM('o036542, 16'o000000);
`MEM('o036544, 16'o000000);
`MEM('o036546, 16'o000000);
`MEM('o036550, 16'o000000);
`MEM('o036552, 16'o000000);
`MEM('o036554, 16'o000000);
`MEM('o036556, 16'o000000);
`MEM('o036560, 16'o000000);
`MEM('o036562, 16'o000000);
`MEM('o036564, 16'o000000);
`MEM('o036566, 16'o000000);
`MEM('o036570, 16'o000000);
`MEM('o036572, 16'o000000);
`MEM('o036574, 16'o000000);
`MEM('o036576, 16'o000000);
`MEM('o036600, 16'o000000);
`MEM('o036602, 16'o000000);
`MEM('o036604, 16'o000000);
`MEM('o036606, 16'o000000);
`MEM('o036610, 16'o000000);
`MEM('o036612, 16'o000000);
`MEM('o036614, 16'o000000);
`MEM('o036616, 16'o000000);
`MEM('o036620, 16'o000000);
`MEM('o036622, 16'o000000);
`MEM('o036624, 16'o000000);
`MEM('o036626, 16'o000000);
`MEM('o036630, 16'o000000);
`MEM('o036632, 16'o000000);
`MEM('o036634, 16'o000000);
`MEM('o036636, 16'o000000);
`MEM('o036640, 16'o000000);
`MEM('o036642, 16'o000000);
`MEM('o036644, 16'o000000);
`MEM('o036646, 16'o000000);
`MEM('o036650, 16'o000000);
`MEM('o036652, 16'o000000);
`MEM('o036654, 16'o000000);
`MEM('o036656, 16'o000000);
`MEM('o036660, 16'o000000);
`MEM('o036662, 16'o000000);
`MEM('o036664, 16'o000000);
`MEM('o036666, 16'o000000);
`MEM('o036670, 16'o000000);
`MEM('o036672, 16'o000000);
`MEM('o036674, 16'o000000);
`MEM('o036676, 16'o000000);
`MEM('o036700, 16'o000000);
`MEM('o036702, 16'o000000);
`MEM('o036704, 16'o000000);
`MEM('o036706, 16'o000000);
`MEM('o036710, 16'o000000);
`MEM('o036712, 16'o000000);
`MEM('o036714, 16'o000000);
`MEM('o036716, 16'o000000);
`MEM('o036720, 16'o000000);
`MEM('o036722, 16'o000000);
`MEM('o036724, 16'o000000);
`MEM('o036726, 16'o000000);
`MEM('o036730, 16'o000000);
`MEM('o036732, 16'o000000);
`MEM('o036734, 16'o000000);
`MEM('o036736, 16'o000000);
`MEM('o036740, 16'o000000);
`MEM('o036742, 16'o000000);
`MEM('o036744, 16'o000000);
`MEM('o036746, 16'o000000);
`MEM('o036750, 16'o000000);
`MEM('o036752, 16'o000000);
`MEM('o036754, 16'o000000);
`MEM('o036756, 16'o000000);
`MEM('o036760, 16'o000000);
`MEM('o036762, 16'o000000);
`MEM('o036764, 16'o000000);
`MEM('o036766, 16'o000000);
`MEM('o036770, 16'o000000);
`MEM('o036772, 16'o000000);
`MEM('o036774, 16'o000000);
`MEM('o036776, 16'o000000);
`MEM('o037000, 16'o000000);
`MEM('o037002, 16'o000000);
`MEM('o037004, 16'o000000);
`MEM('o037006, 16'o000000);
`MEM('o037010, 16'o000000);
`MEM('o037012, 16'o000000);
`MEM('o037014, 16'o000000);
`MEM('o037016, 16'o000000);
`MEM('o037020, 16'o000000);
`MEM('o037022, 16'o000000);
`MEM('o037024, 16'o000000);
`MEM('o037026, 16'o000000);
`MEM('o037030, 16'o000000);
`MEM('o037032, 16'o000000);
`MEM('o037034, 16'o000000);
`MEM('o037036, 16'o000000);
`MEM('o037040, 16'o000000);
`MEM('o037042, 16'o000000);
`MEM('o037044, 16'o000000);
`MEM('o037046, 16'o000000);
`MEM('o037050, 16'o000000);
`MEM('o037052, 16'o000000);
`MEM('o037054, 16'o000000);
`MEM('o037056, 16'o000000);
`MEM('o037060, 16'o000000);
`MEM('o037062, 16'o000000);
`MEM('o037064, 16'o000000);
`MEM('o037066, 16'o000000);
`MEM('o037070, 16'o000000);
`MEM('o037072, 16'o000000);
`MEM('o037074, 16'o000000);
`MEM('o037076, 16'o000000);
`MEM('o037100, 16'o000000);
`MEM('o037102, 16'o000000);
`MEM('o037104, 16'o000000);
`MEM('o037106, 16'o000000);
`MEM('o037110, 16'o000000);
`MEM('o037112, 16'o000000);
`MEM('o037114, 16'o000000);
`MEM('o037116, 16'o000000);
`MEM('o037120, 16'o000000);
`MEM('o037122, 16'o000000);
`MEM('o037124, 16'o000000);
`MEM('o037126, 16'o000000);
`MEM('o037130, 16'o000000);
`MEM('o037132, 16'o000000);
`MEM('o037134, 16'o000000);
`MEM('o037136, 16'o000000);
`MEM('o037140, 16'o000000);
`MEM('o037142, 16'o000000);
`MEM('o037144, 16'o000000);
`MEM('o037146, 16'o000000);
`MEM('o037150, 16'o000000);
`MEM('o037152, 16'o000000);
`MEM('o037154, 16'o000000);
`MEM('o037156, 16'o000000);
`MEM('o037160, 16'o000000);
`MEM('o037162, 16'o000000);
`MEM('o037164, 16'o000000);
`MEM('o037166, 16'o000000);
`MEM('o037170, 16'o000000);
`MEM('o037172, 16'o000000);
`MEM('o037174, 16'o000000);
`MEM('o037176, 16'o000000);
`MEM('o037200, 16'o000000);
`MEM('o037202, 16'o000000);
`MEM('o037204, 16'o000000);
`MEM('o037206, 16'o000000);
`MEM('o037210, 16'o000000);
`MEM('o037212, 16'o000000);
`MEM('o037214, 16'o000000);
`MEM('o037216, 16'o000000);
`MEM('o037220, 16'o000000);
`MEM('o037222, 16'o000000);
`MEM('o037224, 16'o000000);
`MEM('o037226, 16'o000000);
`MEM('o037230, 16'o000000);
`MEM('o037232, 16'o000000);
`MEM('o037234, 16'o000000);
`MEM('o037236, 16'o000000);
`MEM('o037240, 16'o000000);
`MEM('o037242, 16'o000000);
`MEM('o037244, 16'o000000);
`MEM('o037246, 16'o000000);
`MEM('o037250, 16'o000000);
`MEM('o037252, 16'o000000);
`MEM('o037254, 16'o000000);
`MEM('o037256, 16'o000000);
`MEM('o037260, 16'o000000);
`MEM('o037262, 16'o000000);
`MEM('o037264, 16'o000000);
`MEM('o037266, 16'o000000);
`MEM('o037270, 16'o000000);
`MEM('o037272, 16'o000000);
`MEM('o037274, 16'o000000);
`MEM('o037276, 16'o000000);
`MEM('o037300, 16'o000000);
`MEM('o037302, 16'o000000);
`MEM('o037304, 16'o000000);
`MEM('o037306, 16'o000000);
`MEM('o037310, 16'o000000);
`MEM('o037312, 16'o000000);
`MEM('o037314, 16'o000000);
`MEM('o037316, 16'o000000);
`MEM('o037320, 16'o000000);
`MEM('o037322, 16'o000000);
`MEM('o037324, 16'o000000);
`MEM('o037326, 16'o000000);
`MEM('o037330, 16'o000000);
`MEM('o037332, 16'o000000);
`MEM('o037334, 16'o000000);
`MEM('o037336, 16'o000000);
`MEM('o037340, 16'o000000);
`MEM('o037342, 16'o000000);
`MEM('o037344, 16'o000000);
`MEM('o037346, 16'o000000);
`MEM('o037350, 16'o000000);
`MEM('o037352, 16'o000000);
`MEM('o037354, 16'o000000);
`MEM('o037356, 16'o000000);
`MEM('o037360, 16'o000000);
`MEM('o037362, 16'o000000);
`MEM('o037364, 16'o000000);
`MEM('o037366, 16'o000000);
`MEM('o037370, 16'o000000);
`MEM('o037372, 16'o000000);
`MEM('o037374, 16'o000000);
`MEM('o037376, 16'o000000);
`MEM('o037400, 16'o000000);
`MEM('o037402, 16'o000000);
`MEM('o037404, 16'o000000);
`MEM('o037406, 16'o000000);
`MEM('o037410, 16'o000000);
`MEM('o037412, 16'o000000);
`MEM('o037414, 16'o000000);
`MEM('o037416, 16'o000000);
`MEM('o037420, 16'o000000);
`MEM('o037422, 16'o000000);
`MEM('o037424, 16'o000000);
`MEM('o037426, 16'o000000);
`MEM('o037430, 16'o000000);
`MEM('o037432, 16'o000000);
`MEM('o037434, 16'o000000);
`MEM('o037436, 16'o000000);
`MEM('o037440, 16'o000000);
`MEM('o037442, 16'o000000);
`MEM('o037444, 16'o000000);
`MEM('o037446, 16'o000000);
`MEM('o037450, 16'o000000);
`MEM('o037452, 16'o000000);
`MEM('o037454, 16'o000000);
`MEM('o037456, 16'o000000);
`MEM('o037460, 16'o000000);
`MEM('o037462, 16'o000000);
`MEM('o037464, 16'o000000);
`MEM('o037466, 16'o000000);
`MEM('o037470, 16'o000000);
`MEM('o037472, 16'o000000);
`MEM('o037474, 16'o037700);
`MEM('o037476, 16'o000000);
`MEM('o037500, 16'o010706);
`MEM('o037502, 16'o024646);
`MEM('o037504, 16'o010705);
`MEM('o037506, 16'o062705);
`MEM('o037510, 16'o000112);
`MEM('o037512, 16'o005001);
`MEM('o037514, 16'o013716);
`MEM('o037516, 16'o177570);
`MEM('o037520, 16'o006016);
`MEM('o037522, 16'o103402);
`MEM('o037524, 16'o005016);
`MEM('o037526, 16'o000403);
`MEM('o037530, 16'o006316);
`MEM('o037532, 16'o001001);
`MEM('o037534, 16'o010116);
`MEM('o037536, 16'o005000);
`MEM('o037540, 16'o004715);
`MEM('o037542, 16'o105303);
`MEM('o037544, 16'o001374);
`MEM('o037546, 16'o004715);
`MEM('o037550, 16'o004767);
`MEM('o037552, 16'o000074);
`MEM('o037554, 16'o010402);
`MEM('o037556, 16'o162702);
`MEM('o037560, 16'o000004);
`MEM('o037562, 16'o022702);
`MEM('o037564, 16'o000002);
`MEM('o037566, 16'o001441);
`MEM('o037570, 16'o004767);
`MEM('o037572, 16'o000054);
`MEM('o037574, 16'o061604);
`MEM('o037576, 16'o010401);
`MEM('o037600, 16'o004715);
`MEM('o037602, 16'o002004);
`MEM('o037604, 16'o105700);
`MEM('o037606, 16'o001753);
`MEM('o037610, 16'o000000);
`MEM('o037612, 16'o000751);
`MEM('o037614, 16'o110321);
`MEM('o037616, 16'o000770);
`MEM('o037620, 16'o016703);
`MEM('o037622, 16'o000152);
`MEM('o037624, 16'o105213);
`MEM('o037626, 16'o105713);
`MEM('o037630, 16'o100376);
`MEM('o037632, 16'o116303);
`MEM('o037634, 16'o000002);
`MEM('o037636, 16'o060300);
`MEM('o037640, 16'o042703);
`MEM('o037642, 16'o177400);
`MEM('o037644, 16'o005302);
`MEM('o037646, 16'o000207);
`MEM('o037650, 16'o012667);
`MEM('o037652, 16'o000046);
`MEM('o037654, 16'o004715);
`MEM('o037656, 16'o010304);
`MEM('o037660, 16'o004715);
`MEM('o037662, 16'o000303);
`MEM('o037664, 16'o050304);
`MEM('o037666, 16'o016707);
`MEM('o037670, 16'o000030);
`MEM('o037672, 16'o004767);
`MEM('o037674, 16'o177752);
`MEM('o037676, 16'o004715);
`MEM('o037700, 16'o105700);
`MEM('o037702, 16'o001342);
`MEM('o037704, 16'o006204);
`MEM('o037706, 16'o103002);
`MEM('o037710, 16'o000000);
`MEM('o037712, 16'o000700);
`MEM('o037714, 16'o006304);
`MEM('o037716, 16'o061604);
`MEM('o037720, 16'o000114);
`MEM('o037722, 16'o037676);
`MEM('o037724, 16'o012767);
`MEM('o037726, 16'o000352);
`MEM('o037730, 16'o000020);
`MEM('o037732, 16'o012767);
`MEM('o037734, 16'o000765);
`MEM('o037736, 16'o000034);
`MEM('o037740, 16'o000167);
`MEM('o037742, 16'o177532);
`MEM('o037744, 16'o016701);
`MEM('o037746, 16'o000026);
`MEM('o037750, 16'o012702);
`MEM('o037752, 16'o000352);
`MEM('o037754, 16'o005211);
`MEM('o037756, 16'o105711);
`MEM('o037760, 16'o100376);
`MEM('o037762, 16'o116162);
`MEM('o037764, 16'o000002);
`MEM('o037766, 16'o037400);
`MEM('o037770, 16'o005267);
`MEM('o037772, 16'o177756);
`MEM('o037774, 16'o000765);
`MEM('o037776, 16'o177550);
`MEM('o040000, 16'o000000);
`MEM('o040002, 16'o000000);
`MEM('o040004, 16'o000000);
`MEM('o040006, 16'o000000);
`MEM('o040010, 16'o000000);
`MEM('o040012, 16'o000000);
`MEM('o040014, 16'o000000);
`MEM('o040016, 16'o000000);
`MEM('o040020, 16'o000000);
`MEM('o040022, 16'o000000);
`MEM('o040024, 16'o000000);
`MEM('o040026, 16'o000000);
`MEM('o040030, 16'o000000);
`MEM('o040032, 16'o000000);
`MEM('o040034, 16'o000000);
`MEM('o040036, 16'o000000);
`MEM('o040040, 16'o000000);
`MEM('o040042, 16'o000000);
`MEM('o040044, 16'o000000);
`MEM('o040046, 16'o000000);
`MEM('o040050, 16'o000000);
`MEM('o040052, 16'o000000);
`MEM('o040054, 16'o000000);
`MEM('o040056, 16'o000000);
`MEM('o040060, 16'o000000);
`MEM('o040062, 16'o000000);
`MEM('o040064, 16'o000000);
`MEM('o040066, 16'o000000);
`MEM('o040070, 16'o000000);
`MEM('o040072, 16'o000000);
`MEM('o040074, 16'o000000);
`MEM('o040076, 16'o000000);
`MEM('o040100, 16'o000000);
`MEM('o040102, 16'o000000);
`MEM('o040104, 16'o000000);
`MEM('o040106, 16'o000000);
`MEM('o040110, 16'o000000);
`MEM('o040112, 16'o000000);
`MEM('o040114, 16'o000000);
`MEM('o040116, 16'o000000);
`MEM('o040120, 16'o000000);
`MEM('o040122, 16'o000000);
`MEM('o040124, 16'o000000);
`MEM('o040126, 16'o000000);
`MEM('o040130, 16'o000000);
`MEM('o040132, 16'o000000);
`MEM('o040134, 16'o000000);
`MEM('o040136, 16'o000000);
`MEM('o040140, 16'o000000);
`MEM('o040142, 16'o000000);
`MEM('o040144, 16'o000000);
`MEM('o040146, 16'o000000);
`MEM('o040150, 16'o000000);
`MEM('o040152, 16'o000000);
`MEM('o040154, 16'o000000);
`MEM('o040156, 16'o000000);
`MEM('o040160, 16'o000000);
`MEM('o040162, 16'o000000);
`MEM('o040164, 16'o000000);
`MEM('o040166, 16'o000000);
`MEM('o040170, 16'o000000);
`MEM('o040172, 16'o000000);
`MEM('o040174, 16'o000000);
`MEM('o040176, 16'o000000);
`MEM('o040200, 16'o000000);
`MEM('o040202, 16'o000000);
`MEM('o040204, 16'o000000);
`MEM('o040206, 16'o000000);
`MEM('o040210, 16'o000000);
`MEM('o040212, 16'o000000);
`MEM('o040214, 16'o000000);
`MEM('o040216, 16'o000000);
`MEM('o040220, 16'o000000);
`MEM('o040222, 16'o000000);
`MEM('o040224, 16'o000000);
`MEM('o040226, 16'o000000);
`MEM('o040230, 16'o000000);
`MEM('o040232, 16'o000000);
`MEM('o040234, 16'o000000);
`MEM('o040236, 16'o000000);
`MEM('o040240, 16'o000000);
`MEM('o040242, 16'o000000);
`MEM('o040244, 16'o000000);
`MEM('o040246, 16'o000000);
`MEM('o040250, 16'o000000);
`MEM('o040252, 16'o000000);
`MEM('o040254, 16'o000000);
`MEM('o040256, 16'o000000);
`MEM('o040260, 16'o000000);
`MEM('o040262, 16'o000000);
`MEM('o040264, 16'o000000);
`MEM('o040266, 16'o000000);
`MEM('o040270, 16'o000000);
`MEM('o040272, 16'o000000);
`MEM('o040274, 16'o000000);
`MEM('o040276, 16'o000000);
`MEM('o040300, 16'o000000);
`MEM('o040302, 16'o000000);
`MEM('o040304, 16'o000000);
`MEM('o040306, 16'o000000);
`MEM('o040310, 16'o000000);
`MEM('o040312, 16'o000000);
`MEM('o040314, 16'o000000);
`MEM('o040316, 16'o000000);
`MEM('o040320, 16'o000000);
`MEM('o040322, 16'o000000);
`MEM('o040324, 16'o000000);
`MEM('o040326, 16'o000000);
`MEM('o040330, 16'o000000);
`MEM('o040332, 16'o000000);
`MEM('o040334, 16'o000000);
`MEM('o040336, 16'o000000);
`MEM('o040340, 16'o000000);
`MEM('o040342, 16'o000000);
`MEM('o040344, 16'o000000);
`MEM('o040346, 16'o000000);
`MEM('o040350, 16'o000000);
`MEM('o040352, 16'o000000);
`MEM('o040354, 16'o000000);
`MEM('o040356, 16'o000000);
`MEM('o040360, 16'o000000);
`MEM('o040362, 16'o000000);
`MEM('o040364, 16'o000000);
`MEM('o040366, 16'o000000);
`MEM('o040370, 16'o000000);
`MEM('o040372, 16'o000000);
`MEM('o040374, 16'o000000);
`MEM('o040376, 16'o000000);
`MEM('o040400, 16'o000000);
`MEM('o040402, 16'o000000);
`MEM('o040404, 16'o000000);
`MEM('o040406, 16'o000000);
`MEM('o040410, 16'o000000);
`MEM('o040412, 16'o000000);
`MEM('o040414, 16'o000000);
`MEM('o040416, 16'o000000);
`MEM('o040420, 16'o000000);
`MEM('o040422, 16'o000000);
`MEM('o040424, 16'o000000);
`MEM('o040426, 16'o000000);
`MEM('o040430, 16'o000000);
`MEM('o040432, 16'o000000);
`MEM('o040434, 16'o000000);
`MEM('o040436, 16'o000000);
`MEM('o040440, 16'o000000);
`MEM('o040442, 16'o000000);
`MEM('o040444, 16'o000000);
`MEM('o040446, 16'o000000);
`MEM('o040450, 16'o000000);
`MEM('o040452, 16'o000000);
`MEM('o040454, 16'o000000);
`MEM('o040456, 16'o000000);
`MEM('o040460, 16'o000000);
`MEM('o040462, 16'o000000);
`MEM('o040464, 16'o000000);
`MEM('o040466, 16'o000000);
`MEM('o040470, 16'o000000);
`MEM('o040472, 16'o000000);
`MEM('o040474, 16'o000000);
`MEM('o040476, 16'o000000);
`MEM('o040500, 16'o000000);
`MEM('o040502, 16'o000000);
`MEM('o040504, 16'o000000);
`MEM('o040506, 16'o000000);
`MEM('o040510, 16'o000000);
`MEM('o040512, 16'o000000);
`MEM('o040514, 16'o000000);
`MEM('o040516, 16'o000000);
`MEM('o040520, 16'o000000);
`MEM('o040522, 16'o000000);
`MEM('o040524, 16'o000000);
`MEM('o040526, 16'o000000);
`MEM('o040530, 16'o000000);
`MEM('o040532, 16'o000000);
`MEM('o040534, 16'o000000);
`MEM('o040536, 16'o000000);
`MEM('o040540, 16'o000000);
`MEM('o040542, 16'o000000);
`MEM('o040544, 16'o000000);
`MEM('o040546, 16'o000000);
`MEM('o040550, 16'o000000);
`MEM('o040552, 16'o000000);
`MEM('o040554, 16'o000000);
`MEM('o040556, 16'o000000);
`MEM('o040560, 16'o000000);
`MEM('o040562, 16'o000000);
`MEM('o040564, 16'o000000);
`MEM('o040566, 16'o000000);
`MEM('o040570, 16'o000000);
`MEM('o040572, 16'o000000);
`MEM('o040574, 16'o000000);
`MEM('o040576, 16'o000000);
`MEM('o040600, 16'o000000);
`MEM('o040602, 16'o000000);
`MEM('o040604, 16'o000000);
`MEM('o040606, 16'o000000);
`MEM('o040610, 16'o000000);
`MEM('o040612, 16'o000000);
`MEM('o040614, 16'o000000);
`MEM('o040616, 16'o000000);
`MEM('o040620, 16'o000000);
`MEM('o040622, 16'o000000);
`MEM('o040624, 16'o000000);
`MEM('o040626, 16'o000000);
`MEM('o040630, 16'o000000);
`MEM('o040632, 16'o000000);
`MEM('o040634, 16'o000000);
`MEM('o040636, 16'o000000);
`MEM('o040640, 16'o000000);
`MEM('o040642, 16'o000000);
`MEM('o040644, 16'o000000);
`MEM('o040646, 16'o000000);
`MEM('o040650, 16'o000000);
`MEM('o040652, 16'o000000);
`MEM('o040654, 16'o000000);
`MEM('o040656, 16'o000000);
`MEM('o040660, 16'o000000);
`MEM('o040662, 16'o000000);
`MEM('o040664, 16'o000000);
`MEM('o040666, 16'o000000);
`MEM('o040670, 16'o000000);
`MEM('o040672, 16'o000000);
`MEM('o040674, 16'o000000);
`MEM('o040676, 16'o000000);
`MEM('o040700, 16'o000000);
`MEM('o040702, 16'o000000);
`MEM('o040704, 16'o000000);
`MEM('o040706, 16'o000000);
`MEM('o040710, 16'o000000);
`MEM('o040712, 16'o000000);
`MEM('o040714, 16'o000000);
`MEM('o040716, 16'o000000);
`MEM('o040720, 16'o000000);
`MEM('o040722, 16'o000000);
`MEM('o040724, 16'o000000);
`MEM('o040726, 16'o000000);
`MEM('o040730, 16'o000000);
`MEM('o040732, 16'o000000);
`MEM('o040734, 16'o000000);
`MEM('o040736, 16'o000000);
`MEM('o040740, 16'o000000);
`MEM('o040742, 16'o000000);
`MEM('o040744, 16'o000000);
`MEM('o040746, 16'o000000);
`MEM('o040750, 16'o000000);
`MEM('o040752, 16'o000000);
`MEM('o040754, 16'o000000);
`MEM('o040756, 16'o000000);
`MEM('o040760, 16'o000000);
`MEM('o040762, 16'o000000);
`MEM('o040764, 16'o000000);
`MEM('o040766, 16'o000000);
`MEM('o040770, 16'o000000);
`MEM('o040772, 16'o000000);
`MEM('o040774, 16'o000000);
`MEM('o040776, 16'o000000);
`MEM('o041000, 16'o000000);
`MEM('o041002, 16'o000000);
`MEM('o041004, 16'o000000);
`MEM('o041006, 16'o000000);
`MEM('o041010, 16'o000000);
`MEM('o041012, 16'o000000);
`MEM('o041014, 16'o000000);
`MEM('o041016, 16'o000000);
`MEM('o041020, 16'o000000);
`MEM('o041022, 16'o000000);
`MEM('o041024, 16'o000000);
`MEM('o041026, 16'o000000);
`MEM('o041030, 16'o000000);
`MEM('o041032, 16'o000000);
`MEM('o041034, 16'o000000);
`MEM('o041036, 16'o000000);
`MEM('o041040, 16'o000000);
`MEM('o041042, 16'o000000);
`MEM('o041044, 16'o000000);
`MEM('o041046, 16'o000000);
`MEM('o041050, 16'o000000);
`MEM('o041052, 16'o000000);
`MEM('o041054, 16'o000000);
`MEM('o041056, 16'o000000);
`MEM('o041060, 16'o000000);
`MEM('o041062, 16'o000000);
`MEM('o041064, 16'o000000);
`MEM('o041066, 16'o000000);
`MEM('o041070, 16'o000000);
`MEM('o041072, 16'o000000);
`MEM('o041074, 16'o000000);
`MEM('o041076, 16'o000000);
`MEM('o041100, 16'o000000);
`MEM('o041102, 16'o000000);
`MEM('o041104, 16'o000000);
`MEM('o041106, 16'o000000);
`MEM('o041110, 16'o000000);
`MEM('o041112, 16'o000000);
`MEM('o041114, 16'o000000);
`MEM('o041116, 16'o000000);
`MEM('o041120, 16'o000000);
`MEM('o041122, 16'o000000);
`MEM('o041124, 16'o000000);
`MEM('o041126, 16'o000000);
`MEM('o041130, 16'o000000);
`MEM('o041132, 16'o000000);
`MEM('o041134, 16'o000000);
`MEM('o041136, 16'o000000);
`MEM('o041140, 16'o000000);
`MEM('o041142, 16'o000000);
`MEM('o041144, 16'o000000);
`MEM('o041146, 16'o000000);
`MEM('o041150, 16'o000000);
`MEM('o041152, 16'o000000);
`MEM('o041154, 16'o000000);
`MEM('o041156, 16'o000000);
`MEM('o041160, 16'o000000);
`MEM('o041162, 16'o000000);
`MEM('o041164, 16'o000000);
`MEM('o041166, 16'o000000);
`MEM('o041170, 16'o000000);
`MEM('o041172, 16'o000000);
`MEM('o041174, 16'o000000);
`MEM('o041176, 16'o000000);
`MEM('o041200, 16'o000000);
`MEM('o041202, 16'o000000);
`MEM('o041204, 16'o000000);
`MEM('o041206, 16'o000000);
`MEM('o041210, 16'o000000);
`MEM('o041212, 16'o000000);
`MEM('o041214, 16'o000000);
`MEM('o041216, 16'o000000);
`MEM('o041220, 16'o000000);
`MEM('o041222, 16'o000000);
`MEM('o041224, 16'o000000);
`MEM('o041226, 16'o000000);
`MEM('o041230, 16'o000000);
`MEM('o041232, 16'o000000);
`MEM('o041234, 16'o000000);
`MEM('o041236, 16'o000000);
`MEM('o041240, 16'o000000);
`MEM('o041242, 16'o000000);
`MEM('o041244, 16'o000000);
`MEM('o041246, 16'o000000);
`MEM('o041250, 16'o000000);
`MEM('o041252, 16'o000000);
`MEM('o041254, 16'o000000);
`MEM('o041256, 16'o000000);
`MEM('o041260, 16'o000000);
`MEM('o041262, 16'o000000);
`MEM('o041264, 16'o000000);
`MEM('o041266, 16'o000000);
`MEM('o041270, 16'o000000);
`MEM('o041272, 16'o000000);
`MEM('o041274, 16'o000000);
`MEM('o041276, 16'o000000);
`MEM('o041300, 16'o000000);
`MEM('o041302, 16'o000000);
`MEM('o041304, 16'o000000);
`MEM('o041306, 16'o000000);
`MEM('o041310, 16'o000000);
`MEM('o041312, 16'o000000);
`MEM('o041314, 16'o000000);
`MEM('o041316, 16'o000000);
`MEM('o041320, 16'o000000);
`MEM('o041322, 16'o000000);
`MEM('o041324, 16'o000000);
`MEM('o041326, 16'o000000);
`MEM('o041330, 16'o000000);
`MEM('o041332, 16'o000000);
`MEM('o041334, 16'o000000);
`MEM('o041336, 16'o000000);
`MEM('o041340, 16'o000000);
`MEM('o041342, 16'o000000);
`MEM('o041344, 16'o000000);
`MEM('o041346, 16'o000000);
`MEM('o041350, 16'o000000);
`MEM('o041352, 16'o000000);
`MEM('o041354, 16'o000000);
`MEM('o041356, 16'o000000);
`MEM('o041360, 16'o000000);
`MEM('o041362, 16'o000000);
`MEM('o041364, 16'o000000);
`MEM('o041366, 16'o000000);
`MEM('o041370, 16'o000000);
`MEM('o041372, 16'o000000);
`MEM('o041374, 16'o000000);
`MEM('o041376, 16'o000000);
`MEM('o041400, 16'o000000);
`MEM('o041402, 16'o000000);
`MEM('o041404, 16'o000000);
`MEM('o041406, 16'o000000);
`MEM('o041410, 16'o000000);
`MEM('o041412, 16'o000000);
`MEM('o041414, 16'o000000);
`MEM('o041416, 16'o000000);
`MEM('o041420, 16'o000000);
`MEM('o041422, 16'o000000);
`MEM('o041424, 16'o000000);
`MEM('o041426, 16'o000000);
`MEM('o041430, 16'o000000);
`MEM('o041432, 16'o000000);
`MEM('o041434, 16'o000000);
`MEM('o041436, 16'o000000);
`MEM('o041440, 16'o000000);
`MEM('o041442, 16'o000000);
`MEM('o041444, 16'o000000);
`MEM('o041446, 16'o000000);
`MEM('o041450, 16'o000000);
`MEM('o041452, 16'o000000);
`MEM('o041454, 16'o000000);
`MEM('o041456, 16'o000000);
`MEM('o041460, 16'o000000);
`MEM('o041462, 16'o000000);
`MEM('o041464, 16'o000000);
`MEM('o041466, 16'o000000);
`MEM('o041470, 16'o000000);
`MEM('o041472, 16'o000000);
`MEM('o041474, 16'o000000);
`MEM('o041476, 16'o000000);
`MEM('o041500, 16'o000000);
`MEM('o041502, 16'o000000);
`MEM('o041504, 16'o000000);
`MEM('o041506, 16'o000000);
`MEM('o041510, 16'o000000);
`MEM('o041512, 16'o000000);
`MEM('o041514, 16'o000000);
`MEM('o041516, 16'o000000);
`MEM('o041520, 16'o000000);
`MEM('o041522, 16'o000000);
`MEM('o041524, 16'o000000);
`MEM('o041526, 16'o000000);
`MEM('o041530, 16'o000000);
`MEM('o041532, 16'o000000);
`MEM('o041534, 16'o000000);
`MEM('o041536, 16'o000000);
`MEM('o041540, 16'o000000);
`MEM('o041542, 16'o000000);
`MEM('o041544, 16'o000000);
`MEM('o041546, 16'o000000);
`MEM('o041550, 16'o000000);
`MEM('o041552, 16'o000000);
`MEM('o041554, 16'o000000);
`MEM('o041556, 16'o000000);
`MEM('o041560, 16'o000000);
`MEM('o041562, 16'o000000);
`MEM('o041564, 16'o000000);
`MEM('o041566, 16'o000000);
`MEM('o041570, 16'o000000);
`MEM('o041572, 16'o000000);
`MEM('o041574, 16'o000000);
`MEM('o041576, 16'o000000);
`MEM('o041600, 16'o000000);
`MEM('o041602, 16'o000000);
`MEM('o041604, 16'o000000);
`MEM('o041606, 16'o000000);
`MEM('o041610, 16'o000000);
`MEM('o041612, 16'o000000);
`MEM('o041614, 16'o000000);
`MEM('o041616, 16'o000000);
`MEM('o041620, 16'o000000);
`MEM('o041622, 16'o000000);
`MEM('o041624, 16'o000000);
`MEM('o041626, 16'o000000);
`MEM('o041630, 16'o000000);
`MEM('o041632, 16'o000000);
`MEM('o041634, 16'o000000);
`MEM('o041636, 16'o000000);
`MEM('o041640, 16'o000000);
`MEM('o041642, 16'o000000);
`MEM('o041644, 16'o000000);
`MEM('o041646, 16'o000000);
`MEM('o041650, 16'o000000);
`MEM('o041652, 16'o000000);
`MEM('o041654, 16'o000000);
`MEM('o041656, 16'o000000);
`MEM('o041660, 16'o000000);
`MEM('o041662, 16'o000000);
`MEM('o041664, 16'o000000);
`MEM('o041666, 16'o000000);
`MEM('o041670, 16'o000000);
`MEM('o041672, 16'o000000);
`MEM('o041674, 16'o000000);
`MEM('o041676, 16'o000000);
`MEM('o041700, 16'o000000);
`MEM('o041702, 16'o000000);
`MEM('o041704, 16'o000000);
`MEM('o041706, 16'o000000);
`MEM('o041710, 16'o000000);
`MEM('o041712, 16'o000000);
`MEM('o041714, 16'o000000);
`MEM('o041716, 16'o000000);
`MEM('o041720, 16'o000000);
`MEM('o041722, 16'o000000);
`MEM('o041724, 16'o000000);
`MEM('o041726, 16'o000000);
`MEM('o041730, 16'o000000);
`MEM('o041732, 16'o000000);
`MEM('o041734, 16'o000000);
`MEM('o041736, 16'o000000);
`MEM('o041740, 16'o000000);
`MEM('o041742, 16'o000000);
`MEM('o041744, 16'o000000);
`MEM('o041746, 16'o000000);
`MEM('o041750, 16'o000000);
`MEM('o041752, 16'o000000);
`MEM('o041754, 16'o000000);
`MEM('o041756, 16'o000000);
`MEM('o041760, 16'o000000);
`MEM('o041762, 16'o000000);
`MEM('o041764, 16'o000000);
`MEM('o041766, 16'o000000);
`MEM('o041770, 16'o000000);
`MEM('o041772, 16'o000000);
`MEM('o041774, 16'o000000);
`MEM('o041776, 16'o000000);
`MEM('o042000, 16'o000000);
`MEM('o042002, 16'o000000);
`MEM('o042004, 16'o000000);
`MEM('o042006, 16'o000000);
`MEM('o042010, 16'o000000);
`MEM('o042012, 16'o000000);
`MEM('o042014, 16'o000000);
`MEM('o042016, 16'o000000);
`MEM('o042020, 16'o000000);
`MEM('o042022, 16'o000000);
`MEM('o042024, 16'o000000);
`MEM('o042026, 16'o000000);
`MEM('o042030, 16'o000000);
`MEM('o042032, 16'o000000);
`MEM('o042034, 16'o000000);
`MEM('o042036, 16'o000000);
`MEM('o042040, 16'o000000);
`MEM('o042042, 16'o000000);
`MEM('o042044, 16'o000000);
`MEM('o042046, 16'o000000);
`MEM('o042050, 16'o000000);
`MEM('o042052, 16'o000000);
`MEM('o042054, 16'o000000);
`MEM('o042056, 16'o000000);
`MEM('o042060, 16'o000000);
`MEM('o042062, 16'o000000);
`MEM('o042064, 16'o000000);
`MEM('o042066, 16'o000000);
`MEM('o042070, 16'o000000);
`MEM('o042072, 16'o000000);
`MEM('o042074, 16'o000000);
`MEM('o042076, 16'o000000);
`MEM('o042100, 16'o000000);
`MEM('o042102, 16'o000000);
`MEM('o042104, 16'o000000);
`MEM('o042106, 16'o000000);
`MEM('o042110, 16'o000000);
`MEM('o042112, 16'o000000);
`MEM('o042114, 16'o000000);
`MEM('o042116, 16'o000000);
`MEM('o042120, 16'o000000);
`MEM('o042122, 16'o000000);
`MEM('o042124, 16'o000000);
`MEM('o042126, 16'o000000);
`MEM('o042130, 16'o000000);
`MEM('o042132, 16'o000000);
`MEM('o042134, 16'o000000);
`MEM('o042136, 16'o000000);
`MEM('o042140, 16'o000000);
`MEM('o042142, 16'o000000);
`MEM('o042144, 16'o000000);
`MEM('o042146, 16'o000000);
`MEM('o042150, 16'o000000);
`MEM('o042152, 16'o000000);
`MEM('o042154, 16'o000000);
`MEM('o042156, 16'o000000);
`MEM('o042160, 16'o000000);
`MEM('o042162, 16'o000000);
`MEM('o042164, 16'o000000);
`MEM('o042166, 16'o000000);
`MEM('o042170, 16'o000000);
`MEM('o042172, 16'o000000);
`MEM('o042174, 16'o000000);
`MEM('o042176, 16'o000000);
`MEM('o042200, 16'o000000);
`MEM('o042202, 16'o000000);
`MEM('o042204, 16'o000000);
`MEM('o042206, 16'o000000);
`MEM('o042210, 16'o000000);
`MEM('o042212, 16'o000000);
`MEM('o042214, 16'o000000);
`MEM('o042216, 16'o000000);
`MEM('o042220, 16'o000000);
`MEM('o042222, 16'o000000);
`MEM('o042224, 16'o000000);
`MEM('o042226, 16'o000000);
`MEM('o042230, 16'o000000);
`MEM('o042232, 16'o000000);
`MEM('o042234, 16'o000000);
`MEM('o042236, 16'o000000);
`MEM('o042240, 16'o000000);
`MEM('o042242, 16'o000000);
`MEM('o042244, 16'o000000);
`MEM('o042246, 16'o000000);
`MEM('o042250, 16'o000000);
`MEM('o042252, 16'o000000);
`MEM('o042254, 16'o000000);
`MEM('o042256, 16'o000000);
`MEM('o042260, 16'o000000);
`MEM('o042262, 16'o000000);
`MEM('o042264, 16'o000000);
`MEM('o042266, 16'o000000);
`MEM('o042270, 16'o000000);
`MEM('o042272, 16'o000000);
`MEM('o042274, 16'o000000);
`MEM('o042276, 16'o000000);
`MEM('o042300, 16'o000000);
`MEM('o042302, 16'o000000);
`MEM('o042304, 16'o000000);
`MEM('o042306, 16'o000000);
`MEM('o042310, 16'o000000);
`MEM('o042312, 16'o000000);
`MEM('o042314, 16'o000000);
`MEM('o042316, 16'o000000);
`MEM('o042320, 16'o000000);
`MEM('o042322, 16'o000000);
`MEM('o042324, 16'o000000);
`MEM('o042326, 16'o000000);
`MEM('o042330, 16'o000000);
`MEM('o042332, 16'o000000);
`MEM('o042334, 16'o000000);
`MEM('o042336, 16'o000000);
`MEM('o042340, 16'o000000);
`MEM('o042342, 16'o000000);
`MEM('o042344, 16'o000000);
`MEM('o042346, 16'o000000);
`MEM('o042350, 16'o000000);
`MEM('o042352, 16'o000000);
`MEM('o042354, 16'o000000);
`MEM('o042356, 16'o000000);
`MEM('o042360, 16'o000000);
`MEM('o042362, 16'o000000);
`MEM('o042364, 16'o000000);
`MEM('o042366, 16'o000000);
`MEM('o042370, 16'o000000);
`MEM('o042372, 16'o000000);
`MEM('o042374, 16'o000000);
`MEM('o042376, 16'o000000);
`MEM('o042400, 16'o000000);
`MEM('o042402, 16'o000000);
`MEM('o042404, 16'o000000);
`MEM('o042406, 16'o000000);
`MEM('o042410, 16'o000000);
`MEM('o042412, 16'o000000);
`MEM('o042414, 16'o000000);
`MEM('o042416, 16'o000000);
`MEM('o042420, 16'o000000);
`MEM('o042422, 16'o000000);
`MEM('o042424, 16'o000000);
`MEM('o042426, 16'o000000);
`MEM('o042430, 16'o000000);
`MEM('o042432, 16'o000000);
`MEM('o042434, 16'o000000);
`MEM('o042436, 16'o000000);
`MEM('o042440, 16'o000000);
`MEM('o042442, 16'o000000);
`MEM('o042444, 16'o000000);
`MEM('o042446, 16'o000000);
`MEM('o042450, 16'o000000);
`MEM('o042452, 16'o000000);
`MEM('o042454, 16'o000000);
`MEM('o042456, 16'o000000);
`MEM('o042460, 16'o000000);
`MEM('o042462, 16'o000000);
`MEM('o042464, 16'o000000);
`MEM('o042466, 16'o000000);
`MEM('o042470, 16'o000000);
`MEM('o042472, 16'o000000);
`MEM('o042474, 16'o000000);
`MEM('o042476, 16'o000000);
`MEM('o042500, 16'o000000);
`MEM('o042502, 16'o000000);
`MEM('o042504, 16'o000000);
`MEM('o042506, 16'o000000);
`MEM('o042510, 16'o000000);
`MEM('o042512, 16'o000000);
`MEM('o042514, 16'o000000);
`MEM('o042516, 16'o000000);
`MEM('o042520, 16'o000000);
`MEM('o042522, 16'o000000);
`MEM('o042524, 16'o000000);
`MEM('o042526, 16'o000000);
`MEM('o042530, 16'o000000);
`MEM('o042532, 16'o000000);
`MEM('o042534, 16'o000000);
`MEM('o042536, 16'o000000);
`MEM('o042540, 16'o000000);
`MEM('o042542, 16'o000000);
`MEM('o042544, 16'o000000);
`MEM('o042546, 16'o000000);
`MEM('o042550, 16'o000000);
`MEM('o042552, 16'o000000);
`MEM('o042554, 16'o000000);
`MEM('o042556, 16'o000000);
`MEM('o042560, 16'o000000);
`MEM('o042562, 16'o000000);
`MEM('o042564, 16'o000000);
`MEM('o042566, 16'o000000);
`MEM('o042570, 16'o000000);
`MEM('o042572, 16'o000000);
`MEM('o042574, 16'o000000);
`MEM('o042576, 16'o000000);
`MEM('o042600, 16'o000000);
`MEM('o042602, 16'o000000);
`MEM('o042604, 16'o000000);
`MEM('o042606, 16'o000000);
`MEM('o042610, 16'o000000);
`MEM('o042612, 16'o000000);
`MEM('o042614, 16'o000000);
`MEM('o042616, 16'o000000);
`MEM('o042620, 16'o000000);
`MEM('o042622, 16'o000000);
`MEM('o042624, 16'o000000);
`MEM('o042626, 16'o000000);
`MEM('o042630, 16'o000000);
`MEM('o042632, 16'o000000);
`MEM('o042634, 16'o000000);
`MEM('o042636, 16'o000000);
`MEM('o042640, 16'o000000);
`MEM('o042642, 16'o000000);
`MEM('o042644, 16'o000000);
`MEM('o042646, 16'o000000);
`MEM('o042650, 16'o000000);
`MEM('o042652, 16'o000000);
`MEM('o042654, 16'o000000);
`MEM('o042656, 16'o000000);
`MEM('o042660, 16'o000000);
`MEM('o042662, 16'o000000);
`MEM('o042664, 16'o000000);
`MEM('o042666, 16'o000000);
`MEM('o042670, 16'o000000);
`MEM('o042672, 16'o000000);
`MEM('o042674, 16'o000000);
`MEM('o042676, 16'o000000);
`MEM('o042700, 16'o000000);
`MEM('o042702, 16'o000000);
`MEM('o042704, 16'o000000);
`MEM('o042706, 16'o000000);
`MEM('o042710, 16'o000000);
`MEM('o042712, 16'o000000);
`MEM('o042714, 16'o000000);
`MEM('o042716, 16'o000000);
`MEM('o042720, 16'o000000);
`MEM('o042722, 16'o000000);
`MEM('o042724, 16'o000000);
`MEM('o042726, 16'o000000);
`MEM('o042730, 16'o000000);
`MEM('o042732, 16'o000000);
`MEM('o042734, 16'o000000);
`MEM('o042736, 16'o000000);
`MEM('o042740, 16'o000000);
`MEM('o042742, 16'o000000);
`MEM('o042744, 16'o000000);
`MEM('o042746, 16'o000000);
`MEM('o042750, 16'o000000);
`MEM('o042752, 16'o000000);
`MEM('o042754, 16'o000000);
`MEM('o042756, 16'o000000);
`MEM('o042760, 16'o000000);
`MEM('o042762, 16'o000000);
`MEM('o042764, 16'o000000);
`MEM('o042766, 16'o000000);
`MEM('o042770, 16'o000000);
`MEM('o042772, 16'o000000);
`MEM('o042774, 16'o000000);
`MEM('o042776, 16'o000000);
`MEM('o043000, 16'o000000);
`MEM('o043002, 16'o000000);
`MEM('o043004, 16'o000000);
`MEM('o043006, 16'o000000);
`MEM('o043010, 16'o000000);
`MEM('o043012, 16'o000000);
`MEM('o043014, 16'o000000);
`MEM('o043016, 16'o000000);
`MEM('o043020, 16'o000000);
`MEM('o043022, 16'o000000);
`MEM('o043024, 16'o000000);
`MEM('o043026, 16'o000000);
`MEM('o043030, 16'o000000);
`MEM('o043032, 16'o000000);
`MEM('o043034, 16'o000000);
`MEM('o043036, 16'o000000);
`MEM('o043040, 16'o000000);
`MEM('o043042, 16'o000000);
`MEM('o043044, 16'o000000);
`MEM('o043046, 16'o000000);
`MEM('o043050, 16'o000000);
`MEM('o043052, 16'o000000);
`MEM('o043054, 16'o000000);
`MEM('o043056, 16'o000000);
`MEM('o043060, 16'o000000);
`MEM('o043062, 16'o000000);
`MEM('o043064, 16'o000000);
`MEM('o043066, 16'o000000);
`MEM('o043070, 16'o000000);
`MEM('o043072, 16'o000000);
`MEM('o043074, 16'o000000);
`MEM('o043076, 16'o000000);
`MEM('o043100, 16'o000000);
`MEM('o043102, 16'o000000);
`MEM('o043104, 16'o000000);
`MEM('o043106, 16'o000000);
`MEM('o043110, 16'o000000);
`MEM('o043112, 16'o000000);
`MEM('o043114, 16'o000000);
`MEM('o043116, 16'o000000);
`MEM('o043120, 16'o000000);
`MEM('o043122, 16'o000000);
`MEM('o043124, 16'o000000);
`MEM('o043126, 16'o000000);
`MEM('o043130, 16'o000000);
`MEM('o043132, 16'o000000);
`MEM('o043134, 16'o000000);
`MEM('o043136, 16'o000000);
`MEM('o043140, 16'o000000);
`MEM('o043142, 16'o000000);
`MEM('o043144, 16'o000000);
`MEM('o043146, 16'o000000);
`MEM('o043150, 16'o000000);
`MEM('o043152, 16'o000000);
`MEM('o043154, 16'o000000);
`MEM('o043156, 16'o000000);
`MEM('o043160, 16'o000000);
`MEM('o043162, 16'o000000);
`MEM('o043164, 16'o000000);
`MEM('o043166, 16'o000000);
`MEM('o043170, 16'o000000);
`MEM('o043172, 16'o000000);
`MEM('o043174, 16'o000000);
`MEM('o043176, 16'o000000);
`MEM('o043200, 16'o000000);
`MEM('o043202, 16'o000000);
`MEM('o043204, 16'o000000);
`MEM('o043206, 16'o000000);
`MEM('o043210, 16'o000000);
`MEM('o043212, 16'o000000);
`MEM('o043214, 16'o000000);
`MEM('o043216, 16'o000000);
`MEM('o043220, 16'o000000);
`MEM('o043222, 16'o000000);
`MEM('o043224, 16'o000000);
`MEM('o043226, 16'o000000);
`MEM('o043230, 16'o000000);
`MEM('o043232, 16'o000000);
`MEM('o043234, 16'o000000);
`MEM('o043236, 16'o000000);
`MEM('o043240, 16'o000000);
`MEM('o043242, 16'o000000);
`MEM('o043244, 16'o000000);
`MEM('o043246, 16'o000000);
`MEM('o043250, 16'o000000);
`MEM('o043252, 16'o000000);
`MEM('o043254, 16'o000000);
`MEM('o043256, 16'o000000);
`MEM('o043260, 16'o000000);
`MEM('o043262, 16'o000000);
`MEM('o043264, 16'o000000);
`MEM('o043266, 16'o000000);
`MEM('o043270, 16'o000000);
`MEM('o043272, 16'o000000);
`MEM('o043274, 16'o000000);
`MEM('o043276, 16'o000000);
`MEM('o043300, 16'o000000);
`MEM('o043302, 16'o000000);
`MEM('o043304, 16'o000000);
`MEM('o043306, 16'o000000);
`MEM('o043310, 16'o000000);
`MEM('o043312, 16'o000000);
`MEM('o043314, 16'o000000);
`MEM('o043316, 16'o000000);
`MEM('o043320, 16'o000000);
`MEM('o043322, 16'o000000);
`MEM('o043324, 16'o000000);
`MEM('o043326, 16'o000000);
`MEM('o043330, 16'o000000);
`MEM('o043332, 16'o000000);
`MEM('o043334, 16'o000000);
`MEM('o043336, 16'o000000);
`MEM('o043340, 16'o000000);
`MEM('o043342, 16'o000000);
`MEM('o043344, 16'o000000);
`MEM('o043346, 16'o000000);
`MEM('o043350, 16'o000000);
`MEM('o043352, 16'o000000);
`MEM('o043354, 16'o000000);
`MEM('o043356, 16'o000000);
`MEM('o043360, 16'o000000);
`MEM('o043362, 16'o000000);
`MEM('o043364, 16'o000000);
`MEM('o043366, 16'o000000);
`MEM('o043370, 16'o000000);
`MEM('o043372, 16'o000000);
`MEM('o043374, 16'o000000);
`MEM('o043376, 16'o000000);
`MEM('o043400, 16'o000000);
`MEM('o043402, 16'o000000);
`MEM('o043404, 16'o000000);
`MEM('o043406, 16'o000000);
`MEM('o043410, 16'o000000);
`MEM('o043412, 16'o000000);
`MEM('o043414, 16'o000000);
`MEM('o043416, 16'o000000);
`MEM('o043420, 16'o000000);
`MEM('o043422, 16'o000000);
`MEM('o043424, 16'o000000);
`MEM('o043426, 16'o000000);
`MEM('o043430, 16'o000000);
`MEM('o043432, 16'o000000);
`MEM('o043434, 16'o000000);
`MEM('o043436, 16'o000000);
`MEM('o043440, 16'o000000);
`MEM('o043442, 16'o000000);
`MEM('o043444, 16'o000000);
`MEM('o043446, 16'o000000);
`MEM('o043450, 16'o000000);
`MEM('o043452, 16'o000000);
`MEM('o043454, 16'o000000);
`MEM('o043456, 16'o000000);
`MEM('o043460, 16'o000000);
`MEM('o043462, 16'o000000);
`MEM('o043464, 16'o000000);
`MEM('o043466, 16'o000000);
`MEM('o043470, 16'o000000);
`MEM('o043472, 16'o000000);
`MEM('o043474, 16'o000000);
`MEM('o043476, 16'o000000);
`MEM('o043500, 16'o000000);
`MEM('o043502, 16'o000000);
`MEM('o043504, 16'o000000);
`MEM('o043506, 16'o000000);
`MEM('o043510, 16'o000000);
`MEM('o043512, 16'o000000);
`MEM('o043514, 16'o000000);
`MEM('o043516, 16'o000000);
`MEM('o043520, 16'o000000);
`MEM('o043522, 16'o000000);
`MEM('o043524, 16'o000000);
`MEM('o043526, 16'o000000);
`MEM('o043530, 16'o000000);
`MEM('o043532, 16'o000000);
`MEM('o043534, 16'o000000);
`MEM('o043536, 16'o000000);
`MEM('o043540, 16'o000000);
`MEM('o043542, 16'o000000);
`MEM('o043544, 16'o000000);
`MEM('o043546, 16'o000000);
`MEM('o043550, 16'o000000);
`MEM('o043552, 16'o000000);
`MEM('o043554, 16'o000000);
`MEM('o043556, 16'o000000);
`MEM('o043560, 16'o000000);
`MEM('o043562, 16'o000000);
`MEM('o043564, 16'o000000);
`MEM('o043566, 16'o000000);
`MEM('o043570, 16'o000000);
`MEM('o043572, 16'o000000);
`MEM('o043574, 16'o000000);
`MEM('o043576, 16'o000000);
`MEM('o043600, 16'o000000);
`MEM('o043602, 16'o000000);
`MEM('o043604, 16'o000000);
`MEM('o043606, 16'o000000);
`MEM('o043610, 16'o000000);
`MEM('o043612, 16'o000000);
`MEM('o043614, 16'o000000);
`MEM('o043616, 16'o000000);
`MEM('o043620, 16'o000000);
`MEM('o043622, 16'o000000);
`MEM('o043624, 16'o000000);
`MEM('o043626, 16'o000000);
`MEM('o043630, 16'o000000);
`MEM('o043632, 16'o000000);
`MEM('o043634, 16'o000000);
`MEM('o043636, 16'o000000);
`MEM('o043640, 16'o000000);
`MEM('o043642, 16'o000000);
`MEM('o043644, 16'o000000);
`MEM('o043646, 16'o000000);
`MEM('o043650, 16'o000000);
`MEM('o043652, 16'o000000);
`MEM('o043654, 16'o000000);
`MEM('o043656, 16'o000000);
`MEM('o043660, 16'o000000);
`MEM('o043662, 16'o000000);
`MEM('o043664, 16'o000000);
`MEM('o043666, 16'o000000);
`MEM('o043670, 16'o000000);
`MEM('o043672, 16'o000000);
`MEM('o043674, 16'o000000);
`MEM('o043676, 16'o000000);
`MEM('o043700, 16'o000000);
`MEM('o043702, 16'o000000);
`MEM('o043704, 16'o000000);
`MEM('o043706, 16'o000000);
`MEM('o043710, 16'o000000);
`MEM('o043712, 16'o000000);
`MEM('o043714, 16'o000000);
`MEM('o043716, 16'o000000);
`MEM('o043720, 16'o000000);
`MEM('o043722, 16'o000000);
`MEM('o043724, 16'o000000);
`MEM('o043726, 16'o000000);
`MEM('o043730, 16'o000000);
`MEM('o043732, 16'o000000);
`MEM('o043734, 16'o000000);
`MEM('o043736, 16'o000000);
`MEM('o043740, 16'o000000);
`MEM('o043742, 16'o000000);
`MEM('o043744, 16'o000000);
`MEM('o043746, 16'o000000);
`MEM('o043750, 16'o000000);
`MEM('o043752, 16'o000000);
`MEM('o043754, 16'o000000);
`MEM('o043756, 16'o000000);
`MEM('o043760, 16'o000000);
`MEM('o043762, 16'o000000);
`MEM('o043764, 16'o000000);
`MEM('o043766, 16'o000000);
`MEM('o043770, 16'o000000);
`MEM('o043772, 16'o000000);
`MEM('o043774, 16'o000000);
`MEM('o043776, 16'o000000);
`MEM('o044000, 16'o000000);
`MEM('o044002, 16'o000000);
`MEM('o044004, 16'o000000);
`MEM('o044006, 16'o000000);
`MEM('o044010, 16'o000000);
`MEM('o044012, 16'o000000);
`MEM('o044014, 16'o000000);
`MEM('o044016, 16'o000000);
`MEM('o044020, 16'o000000);
`MEM('o044022, 16'o000000);
`MEM('o044024, 16'o000000);
`MEM('o044026, 16'o000000);
`MEM('o044030, 16'o000000);
`MEM('o044032, 16'o000000);
`MEM('o044034, 16'o000000);
`MEM('o044036, 16'o000000);
`MEM('o044040, 16'o000000);
`MEM('o044042, 16'o000000);
`MEM('o044044, 16'o000000);
`MEM('o044046, 16'o000000);
`MEM('o044050, 16'o000000);
`MEM('o044052, 16'o000000);
`MEM('o044054, 16'o000000);
`MEM('o044056, 16'o000000);
`MEM('o044060, 16'o000000);
`MEM('o044062, 16'o000000);
`MEM('o044064, 16'o000000);
`MEM('o044066, 16'o000000);
`MEM('o044070, 16'o000000);
`MEM('o044072, 16'o000000);
`MEM('o044074, 16'o000000);
`MEM('o044076, 16'o000000);
`MEM('o044100, 16'o000000);
`MEM('o044102, 16'o000000);
`MEM('o044104, 16'o000000);
`MEM('o044106, 16'o000000);
`MEM('o044110, 16'o000000);
`MEM('o044112, 16'o000000);
`MEM('o044114, 16'o000000);
`MEM('o044116, 16'o000000);
`MEM('o044120, 16'o000000);
`MEM('o044122, 16'o000000);
`MEM('o044124, 16'o000000);
`MEM('o044126, 16'o000000);
`MEM('o044130, 16'o000000);
`MEM('o044132, 16'o000000);
`MEM('o044134, 16'o000000);
`MEM('o044136, 16'o000000);
`MEM('o044140, 16'o000000);
`MEM('o044142, 16'o000000);
`MEM('o044144, 16'o000000);
`MEM('o044146, 16'o000000);
`MEM('o044150, 16'o000000);
`MEM('o044152, 16'o000000);
`MEM('o044154, 16'o000000);
`MEM('o044156, 16'o000000);
`MEM('o044160, 16'o000000);
`MEM('o044162, 16'o000000);
`MEM('o044164, 16'o000000);
`MEM('o044166, 16'o000000);
`MEM('o044170, 16'o000000);
`MEM('o044172, 16'o000000);
`MEM('o044174, 16'o000000);
`MEM('o044176, 16'o000000);
`MEM('o044200, 16'o000000);
`MEM('o044202, 16'o000000);
`MEM('o044204, 16'o000000);
`MEM('o044206, 16'o000000);
`MEM('o044210, 16'o000000);
`MEM('o044212, 16'o000000);
`MEM('o044214, 16'o000000);
`MEM('o044216, 16'o000000);
`MEM('o044220, 16'o000000);
`MEM('o044222, 16'o000000);
`MEM('o044224, 16'o000000);
`MEM('o044226, 16'o000000);
`MEM('o044230, 16'o000000);
`MEM('o044232, 16'o000000);
`MEM('o044234, 16'o000000);
`MEM('o044236, 16'o000000);
`MEM('o044240, 16'o000000);
`MEM('o044242, 16'o000000);
`MEM('o044244, 16'o000000);
`MEM('o044246, 16'o000000);
`MEM('o044250, 16'o000000);
`MEM('o044252, 16'o000000);
`MEM('o044254, 16'o000000);
`MEM('o044256, 16'o000000);
`MEM('o044260, 16'o000000);
`MEM('o044262, 16'o000000);
`MEM('o044264, 16'o000000);
`MEM('o044266, 16'o000000);
`MEM('o044270, 16'o000000);
`MEM('o044272, 16'o000000);
`MEM('o044274, 16'o000000);
`MEM('o044276, 16'o000000);
`MEM('o044300, 16'o000000);
`MEM('o044302, 16'o000000);
`MEM('o044304, 16'o000000);
`MEM('o044306, 16'o000000);
`MEM('o044310, 16'o000000);
`MEM('o044312, 16'o000000);
`MEM('o044314, 16'o000000);
`MEM('o044316, 16'o000000);
`MEM('o044320, 16'o000000);
`MEM('o044322, 16'o000000);
`MEM('o044324, 16'o000000);
`MEM('o044326, 16'o000000);
`MEM('o044330, 16'o000000);
`MEM('o044332, 16'o000000);
`MEM('o044334, 16'o000000);
`MEM('o044336, 16'o000000);
`MEM('o044340, 16'o000000);
`MEM('o044342, 16'o000000);
`MEM('o044344, 16'o000000);
`MEM('o044346, 16'o000000);
`MEM('o044350, 16'o000000);
`MEM('o044352, 16'o000000);
`MEM('o044354, 16'o000000);
`MEM('o044356, 16'o000000);
`MEM('o044360, 16'o000000);
`MEM('o044362, 16'o000000);
`MEM('o044364, 16'o000000);
`MEM('o044366, 16'o000000);
`MEM('o044370, 16'o000000);
`MEM('o044372, 16'o000000);
`MEM('o044374, 16'o000000);
`MEM('o044376, 16'o000000);
`MEM('o044400, 16'o000000);
`MEM('o044402, 16'o000000);
`MEM('o044404, 16'o000000);
`MEM('o044406, 16'o000000);
`MEM('o044410, 16'o000000);
`MEM('o044412, 16'o000000);
`MEM('o044414, 16'o000000);
`MEM('o044416, 16'o000000);
`MEM('o044420, 16'o000000);
`MEM('o044422, 16'o000000);
`MEM('o044424, 16'o000000);
`MEM('o044426, 16'o000000);
`MEM('o044430, 16'o000000);
`MEM('o044432, 16'o000000);
`MEM('o044434, 16'o000000);
`MEM('o044436, 16'o000000);
`MEM('o044440, 16'o000000);
`MEM('o044442, 16'o000000);
`MEM('o044444, 16'o000000);
`MEM('o044446, 16'o000000);
`MEM('o044450, 16'o000000);
`MEM('o044452, 16'o000000);
`MEM('o044454, 16'o000000);
`MEM('o044456, 16'o000000);
`MEM('o044460, 16'o000000);
`MEM('o044462, 16'o000000);
`MEM('o044464, 16'o000000);
`MEM('o044466, 16'o000000);
`MEM('o044470, 16'o000000);
`MEM('o044472, 16'o000000);
`MEM('o044474, 16'o000000);
`MEM('o044476, 16'o000000);
`MEM('o044500, 16'o000000);
`MEM('o044502, 16'o000000);
`MEM('o044504, 16'o000000);
`MEM('o044506, 16'o000000);
`MEM('o044510, 16'o000000);
`MEM('o044512, 16'o000000);
`MEM('o044514, 16'o000000);
`MEM('o044516, 16'o000000);
`MEM('o044520, 16'o000000);
`MEM('o044522, 16'o000000);
`MEM('o044524, 16'o000000);
`MEM('o044526, 16'o000000);
`MEM('o044530, 16'o000000);
`MEM('o044532, 16'o000000);
`MEM('o044534, 16'o000000);
`MEM('o044536, 16'o000000);
`MEM('o044540, 16'o000000);
`MEM('o044542, 16'o000000);
`MEM('o044544, 16'o000000);
`MEM('o044546, 16'o000000);
`MEM('o044550, 16'o000000);
`MEM('o044552, 16'o000000);
`MEM('o044554, 16'o000000);
`MEM('o044556, 16'o000000);
`MEM('o044560, 16'o000000);
`MEM('o044562, 16'o000000);
`MEM('o044564, 16'o000000);
`MEM('o044566, 16'o000000);
`MEM('o044570, 16'o000000);
`MEM('o044572, 16'o000000);
`MEM('o044574, 16'o000000);
`MEM('o044576, 16'o000000);
`MEM('o044600, 16'o000000);
`MEM('o044602, 16'o000000);
`MEM('o044604, 16'o000000);
`MEM('o044606, 16'o000000);
`MEM('o044610, 16'o000000);
`MEM('o044612, 16'o000000);
`MEM('o044614, 16'o000000);
`MEM('o044616, 16'o000000);
`MEM('o044620, 16'o000000);
`MEM('o044622, 16'o000000);
`MEM('o044624, 16'o000000);
`MEM('o044626, 16'o000000);
`MEM('o044630, 16'o000000);
`MEM('o044632, 16'o000000);
`MEM('o044634, 16'o000000);
`MEM('o044636, 16'o000000);
`MEM('o044640, 16'o000000);
`MEM('o044642, 16'o000000);
`MEM('o044644, 16'o000000);
`MEM('o044646, 16'o000000);
`MEM('o044650, 16'o000000);
`MEM('o044652, 16'o000000);
`MEM('o044654, 16'o000000);
`MEM('o044656, 16'o000000);
`MEM('o044660, 16'o000000);
`MEM('o044662, 16'o000000);
`MEM('o044664, 16'o000000);
`MEM('o044666, 16'o000000);
`MEM('o044670, 16'o000000);
`MEM('o044672, 16'o000000);
`MEM('o044674, 16'o000000);
`MEM('o044676, 16'o000000);
`MEM('o044700, 16'o000000);
`MEM('o044702, 16'o000000);
`MEM('o044704, 16'o000000);
`MEM('o044706, 16'o000000);
`MEM('o044710, 16'o000000);
`MEM('o044712, 16'o000000);
`MEM('o044714, 16'o000000);
`MEM('o044716, 16'o000000);
`MEM('o044720, 16'o000000);
`MEM('o044722, 16'o000000);
`MEM('o044724, 16'o000000);
`MEM('o044726, 16'o000000);
`MEM('o044730, 16'o000000);
`MEM('o044732, 16'o000000);
`MEM('o044734, 16'o000000);
`MEM('o044736, 16'o000000);
`MEM('o044740, 16'o000000);
`MEM('o044742, 16'o000000);
`MEM('o044744, 16'o000000);
`MEM('o044746, 16'o000000);
`MEM('o044750, 16'o000000);
`MEM('o044752, 16'o000000);
`MEM('o044754, 16'o000000);
`MEM('o044756, 16'o000000);
`MEM('o044760, 16'o000000);
`MEM('o044762, 16'o000000);
`MEM('o044764, 16'o000000);
`MEM('o044766, 16'o000000);
`MEM('o044770, 16'o000000);
`MEM('o044772, 16'o000000);
`MEM('o044774, 16'o000000);
`MEM('o044776, 16'o000000);
`MEM('o045000, 16'o000000);
`MEM('o045002, 16'o000000);
`MEM('o045004, 16'o000000);
`MEM('o045006, 16'o000000);
`MEM('o045010, 16'o000000);
`MEM('o045012, 16'o000000);
`MEM('o045014, 16'o000000);
`MEM('o045016, 16'o000000);
`MEM('o045020, 16'o000000);
`MEM('o045022, 16'o000000);
`MEM('o045024, 16'o000000);
`MEM('o045026, 16'o000000);
`MEM('o045030, 16'o000000);
`MEM('o045032, 16'o000000);
`MEM('o045034, 16'o000000);
`MEM('o045036, 16'o000000);
`MEM('o045040, 16'o000000);
`MEM('o045042, 16'o000000);
`MEM('o045044, 16'o000000);
`MEM('o045046, 16'o000000);
`MEM('o045050, 16'o000000);
`MEM('o045052, 16'o000000);
`MEM('o045054, 16'o000000);
`MEM('o045056, 16'o000000);
`MEM('o045060, 16'o000000);
`MEM('o045062, 16'o000000);
`MEM('o045064, 16'o000000);
`MEM('o045066, 16'o000000);
`MEM('o045070, 16'o000000);
`MEM('o045072, 16'o000000);
`MEM('o045074, 16'o000000);
`MEM('o045076, 16'o000000);
`MEM('o045100, 16'o000000);
`MEM('o045102, 16'o000000);
`MEM('o045104, 16'o000000);
`MEM('o045106, 16'o000000);
`MEM('o045110, 16'o000000);
`MEM('o045112, 16'o000000);
`MEM('o045114, 16'o000000);
`MEM('o045116, 16'o000000);
`MEM('o045120, 16'o000000);
`MEM('o045122, 16'o000000);
`MEM('o045124, 16'o000000);
`MEM('o045126, 16'o000000);
`MEM('o045130, 16'o000000);
`MEM('o045132, 16'o000000);
`MEM('o045134, 16'o000000);
`MEM('o045136, 16'o000000);
`MEM('o045140, 16'o000000);
`MEM('o045142, 16'o000000);
`MEM('o045144, 16'o000000);
`MEM('o045146, 16'o000000);
`MEM('o045150, 16'o000000);
`MEM('o045152, 16'o000000);
`MEM('o045154, 16'o000000);
`MEM('o045156, 16'o000000);
`MEM('o045160, 16'o000000);
`MEM('o045162, 16'o000000);
`MEM('o045164, 16'o000000);
`MEM('o045166, 16'o000000);
`MEM('o045170, 16'o000000);
`MEM('o045172, 16'o000000);
`MEM('o045174, 16'o000000);
`MEM('o045176, 16'o000000);
`MEM('o045200, 16'o000000);
`MEM('o045202, 16'o000000);
`MEM('o045204, 16'o000000);
`MEM('o045206, 16'o000000);
`MEM('o045210, 16'o000000);
`MEM('o045212, 16'o000000);
`MEM('o045214, 16'o000000);
`MEM('o045216, 16'o000000);
`MEM('o045220, 16'o000000);
`MEM('o045222, 16'o000000);
`MEM('o045224, 16'o000000);
`MEM('o045226, 16'o000000);
`MEM('o045230, 16'o000000);
`MEM('o045232, 16'o000000);
`MEM('o045234, 16'o000000);
`MEM('o045236, 16'o000000);
`MEM('o045240, 16'o000000);
`MEM('o045242, 16'o000000);
`MEM('o045244, 16'o000000);
`MEM('o045246, 16'o000000);
`MEM('o045250, 16'o000000);
`MEM('o045252, 16'o000000);
`MEM('o045254, 16'o000000);
`MEM('o045256, 16'o000000);
`MEM('o045260, 16'o000000);
`MEM('o045262, 16'o000000);
`MEM('o045264, 16'o000000);
`MEM('o045266, 16'o000000);
`MEM('o045270, 16'o000000);
`MEM('o045272, 16'o000000);
`MEM('o045274, 16'o000000);
`MEM('o045276, 16'o000000);
`MEM('o045300, 16'o000000);
`MEM('o045302, 16'o000000);
`MEM('o045304, 16'o000000);
`MEM('o045306, 16'o000000);
`MEM('o045310, 16'o000000);
`MEM('o045312, 16'o000000);
`MEM('o045314, 16'o000000);
`MEM('o045316, 16'o000000);
`MEM('o045320, 16'o000000);
`MEM('o045322, 16'o000000);
`MEM('o045324, 16'o000000);
`MEM('o045326, 16'o000000);
`MEM('o045330, 16'o000000);
`MEM('o045332, 16'o000000);
`MEM('o045334, 16'o000000);
`MEM('o045336, 16'o000000);
`MEM('o045340, 16'o000000);
`MEM('o045342, 16'o000000);
`MEM('o045344, 16'o000000);
`MEM('o045346, 16'o000000);
`MEM('o045350, 16'o000000);
`MEM('o045352, 16'o000000);
`MEM('o045354, 16'o000000);
`MEM('o045356, 16'o000000);
`MEM('o045360, 16'o000000);
`MEM('o045362, 16'o000000);
`MEM('o045364, 16'o000000);
`MEM('o045366, 16'o000000);
`MEM('o045370, 16'o000000);
`MEM('o045372, 16'o000000);
`MEM('o045374, 16'o000000);
`MEM('o045376, 16'o000000);
`MEM('o045400, 16'o000000);
`MEM('o045402, 16'o000000);
`MEM('o045404, 16'o000000);
`MEM('o045406, 16'o000000);
`MEM('o045410, 16'o000000);
`MEM('o045412, 16'o000000);
`MEM('o045414, 16'o000000);
`MEM('o045416, 16'o000000);
`MEM('o045420, 16'o000000);
`MEM('o045422, 16'o000000);
`MEM('o045424, 16'o000000);
`MEM('o045426, 16'o000000);
`MEM('o045430, 16'o000000);
`MEM('o045432, 16'o000000);
`MEM('o045434, 16'o000000);
`MEM('o045436, 16'o000000);
`MEM('o045440, 16'o000000);
`MEM('o045442, 16'o000000);
`MEM('o045444, 16'o000000);
`MEM('o045446, 16'o000000);
`MEM('o045450, 16'o000000);
`MEM('o045452, 16'o000000);
`MEM('o045454, 16'o000000);
`MEM('o045456, 16'o000000);
`MEM('o045460, 16'o000000);
`MEM('o045462, 16'o000000);
`MEM('o045464, 16'o000000);
`MEM('o045466, 16'o000000);
`MEM('o045470, 16'o000000);
`MEM('o045472, 16'o000000);
`MEM('o045474, 16'o000000);
`MEM('o045476, 16'o000000);
`MEM('o045500, 16'o000000);
`MEM('o045502, 16'o000000);
`MEM('o045504, 16'o000000);
`MEM('o045506, 16'o000000);
`MEM('o045510, 16'o000000);
`MEM('o045512, 16'o000000);
`MEM('o045514, 16'o000000);
`MEM('o045516, 16'o000000);
`MEM('o045520, 16'o000000);
`MEM('o045522, 16'o000000);
`MEM('o045524, 16'o000000);
`MEM('o045526, 16'o000000);
`MEM('o045530, 16'o000000);
`MEM('o045532, 16'o000000);
`MEM('o045534, 16'o000000);
`MEM('o045536, 16'o000000);
`MEM('o045540, 16'o000000);
`MEM('o045542, 16'o000000);
`MEM('o045544, 16'o000000);
`MEM('o045546, 16'o000000);
`MEM('o045550, 16'o000000);
`MEM('o045552, 16'o000000);
`MEM('o045554, 16'o000000);
`MEM('o045556, 16'o000000);
`MEM('o045560, 16'o000000);
`MEM('o045562, 16'o000000);
`MEM('o045564, 16'o000000);
`MEM('o045566, 16'o000000);
`MEM('o045570, 16'o000000);
`MEM('o045572, 16'o000000);
`MEM('o045574, 16'o000000);
`MEM('o045576, 16'o000000);
`MEM('o045600, 16'o000000);
`MEM('o045602, 16'o000000);
`MEM('o045604, 16'o000000);
`MEM('o045606, 16'o000000);
`MEM('o045610, 16'o000000);
`MEM('o045612, 16'o000000);
`MEM('o045614, 16'o000000);
`MEM('o045616, 16'o000000);
`MEM('o045620, 16'o000000);
`MEM('o045622, 16'o000000);
`MEM('o045624, 16'o000000);
`MEM('o045626, 16'o000000);
`MEM('o045630, 16'o000000);
`MEM('o045632, 16'o000000);
`MEM('o045634, 16'o000000);
`MEM('o045636, 16'o000000);
`MEM('o045640, 16'o000000);
`MEM('o045642, 16'o000000);
`MEM('o045644, 16'o000000);
`MEM('o045646, 16'o000000);
`MEM('o045650, 16'o000000);
`MEM('o045652, 16'o000000);
`MEM('o045654, 16'o000000);
`MEM('o045656, 16'o000000);
`MEM('o045660, 16'o000000);
`MEM('o045662, 16'o000000);
`MEM('o045664, 16'o000000);
`MEM('o045666, 16'o000000);
`MEM('o045670, 16'o000000);
`MEM('o045672, 16'o000000);
`MEM('o045674, 16'o000000);
`MEM('o045676, 16'o000000);
`MEM('o045700, 16'o000000);
`MEM('o045702, 16'o000000);
`MEM('o045704, 16'o000000);
`MEM('o045706, 16'o000000);
`MEM('o045710, 16'o000000);
`MEM('o045712, 16'o000000);
`MEM('o045714, 16'o000000);
`MEM('o045716, 16'o000000);
`MEM('o045720, 16'o000000);
`MEM('o045722, 16'o000000);
`MEM('o045724, 16'o000000);
`MEM('o045726, 16'o000000);
`MEM('o045730, 16'o000000);
`MEM('o045732, 16'o000000);
`MEM('o045734, 16'o000000);
`MEM('o045736, 16'o000000);
`MEM('o045740, 16'o000000);
`MEM('o045742, 16'o000000);
`MEM('o045744, 16'o000000);
`MEM('o045746, 16'o000000);
`MEM('o045750, 16'o000000);
`MEM('o045752, 16'o000000);
`MEM('o045754, 16'o000000);
`MEM('o045756, 16'o000000);
`MEM('o045760, 16'o000000);
`MEM('o045762, 16'o000000);
`MEM('o045764, 16'o000000);
`MEM('o045766, 16'o000000);
`MEM('o045770, 16'o000000);
`MEM('o045772, 16'o000000);
`MEM('o045774, 16'o000000);
`MEM('o045776, 16'o000000);
`MEM('o046000, 16'o000000);
`MEM('o046002, 16'o000000);
`MEM('o046004, 16'o000000);
`MEM('o046006, 16'o000000);
`MEM('o046010, 16'o000000);
`MEM('o046012, 16'o000000);
`MEM('o046014, 16'o000000);
`MEM('o046016, 16'o000000);
`MEM('o046020, 16'o000000);
`MEM('o046022, 16'o000000);
`MEM('o046024, 16'o000000);
`MEM('o046026, 16'o000000);
`MEM('o046030, 16'o000000);
`MEM('o046032, 16'o000000);
`MEM('o046034, 16'o000000);
`MEM('o046036, 16'o000000);
`MEM('o046040, 16'o000000);
`MEM('o046042, 16'o000000);
`MEM('o046044, 16'o000000);
`MEM('o046046, 16'o000000);
`MEM('o046050, 16'o000000);
`MEM('o046052, 16'o000000);
`MEM('o046054, 16'o000000);
`MEM('o046056, 16'o000000);
`MEM('o046060, 16'o000000);
`MEM('o046062, 16'o000000);
`MEM('o046064, 16'o000000);
`MEM('o046066, 16'o000000);
`MEM('o046070, 16'o000000);
`MEM('o046072, 16'o000000);
`MEM('o046074, 16'o000000);
`MEM('o046076, 16'o000000);
`MEM('o046100, 16'o000000);
`MEM('o046102, 16'o000000);
`MEM('o046104, 16'o000000);
`MEM('o046106, 16'o000000);
`MEM('o046110, 16'o000000);
`MEM('o046112, 16'o000000);
`MEM('o046114, 16'o000000);
`MEM('o046116, 16'o000000);
`MEM('o046120, 16'o000000);
`MEM('o046122, 16'o000000);
`MEM('o046124, 16'o000000);
`MEM('o046126, 16'o000000);
`MEM('o046130, 16'o000000);
`MEM('o046132, 16'o000000);
`MEM('o046134, 16'o000000);
`MEM('o046136, 16'o000000);
`MEM('o046140, 16'o000000);
`MEM('o046142, 16'o000000);
`MEM('o046144, 16'o000000);
`MEM('o046146, 16'o000000);
`MEM('o046150, 16'o000000);
`MEM('o046152, 16'o000000);
`MEM('o046154, 16'o000000);
`MEM('o046156, 16'o000000);
`MEM('o046160, 16'o000000);
`MEM('o046162, 16'o000000);
`MEM('o046164, 16'o000000);
`MEM('o046166, 16'o000000);
`MEM('o046170, 16'o000000);
`MEM('o046172, 16'o000000);
`MEM('o046174, 16'o000000);
`MEM('o046176, 16'o000000);
`MEM('o046200, 16'o000000);
`MEM('o046202, 16'o000000);
`MEM('o046204, 16'o000000);
`MEM('o046206, 16'o000000);
`MEM('o046210, 16'o000000);
`MEM('o046212, 16'o000000);
`MEM('o046214, 16'o000000);
`MEM('o046216, 16'o000000);
`MEM('o046220, 16'o000000);
`MEM('o046222, 16'o000000);
`MEM('o046224, 16'o000000);
`MEM('o046226, 16'o000000);
`MEM('o046230, 16'o000000);
`MEM('o046232, 16'o000000);
`MEM('o046234, 16'o000000);
`MEM('o046236, 16'o000000);
`MEM('o046240, 16'o000000);
`MEM('o046242, 16'o000000);
`MEM('o046244, 16'o000000);
`MEM('o046246, 16'o000000);
`MEM('o046250, 16'o000000);
`MEM('o046252, 16'o000000);
`MEM('o046254, 16'o000000);
`MEM('o046256, 16'o000000);
`MEM('o046260, 16'o000000);
`MEM('o046262, 16'o000000);
`MEM('o046264, 16'o000000);
`MEM('o046266, 16'o000000);
`MEM('o046270, 16'o000000);
`MEM('o046272, 16'o000000);
`MEM('o046274, 16'o000000);
`MEM('o046276, 16'o000000);
`MEM('o046300, 16'o000000);
`MEM('o046302, 16'o000000);
`MEM('o046304, 16'o000000);
`MEM('o046306, 16'o000000);
`MEM('o046310, 16'o000000);
`MEM('o046312, 16'o000000);
`MEM('o046314, 16'o000000);
`MEM('o046316, 16'o000000);
`MEM('o046320, 16'o000000);
`MEM('o046322, 16'o000000);
`MEM('o046324, 16'o000000);
`MEM('o046326, 16'o000000);
`MEM('o046330, 16'o000000);
`MEM('o046332, 16'o000000);
`MEM('o046334, 16'o000000);
`MEM('o046336, 16'o000000);
`MEM('o046340, 16'o000000);
`MEM('o046342, 16'o000000);
`MEM('o046344, 16'o000000);
`MEM('o046346, 16'o000000);
`MEM('o046350, 16'o000000);
`MEM('o046352, 16'o000000);
`MEM('o046354, 16'o000000);
`MEM('o046356, 16'o000000);
`MEM('o046360, 16'o000000);
`MEM('o046362, 16'o000000);
`MEM('o046364, 16'o000000);
`MEM('o046366, 16'o000000);
`MEM('o046370, 16'o000000);
`MEM('o046372, 16'o000000);
`MEM('o046374, 16'o000000);
`MEM('o046376, 16'o000000);
`MEM('o046400, 16'o000000);
`MEM('o046402, 16'o000000);
`MEM('o046404, 16'o000000);
`MEM('o046406, 16'o000000);
`MEM('o046410, 16'o000000);
`MEM('o046412, 16'o000000);
`MEM('o046414, 16'o000000);
`MEM('o046416, 16'o000000);
`MEM('o046420, 16'o000000);
`MEM('o046422, 16'o000000);
`MEM('o046424, 16'o000000);
`MEM('o046426, 16'o000000);
`MEM('o046430, 16'o000000);
`MEM('o046432, 16'o000000);
`MEM('o046434, 16'o000000);
`MEM('o046436, 16'o000000);
`MEM('o046440, 16'o000000);
`MEM('o046442, 16'o000000);
`MEM('o046444, 16'o000000);
`MEM('o046446, 16'o000000);
`MEM('o046450, 16'o000000);
`MEM('o046452, 16'o000000);
`MEM('o046454, 16'o000000);
`MEM('o046456, 16'o000000);
`MEM('o046460, 16'o000000);
`MEM('o046462, 16'o000000);
`MEM('o046464, 16'o000000);
`MEM('o046466, 16'o000000);
`MEM('o046470, 16'o000000);
`MEM('o046472, 16'o000000);
`MEM('o046474, 16'o000000);
`MEM('o046476, 16'o000000);
`MEM('o046500, 16'o000000);
`MEM('o046502, 16'o000000);
`MEM('o046504, 16'o000000);
`MEM('o046506, 16'o000000);
`MEM('o046510, 16'o000000);
`MEM('o046512, 16'o000000);
`MEM('o046514, 16'o000000);
`MEM('o046516, 16'o000000);
`MEM('o046520, 16'o000000);
`MEM('o046522, 16'o000000);
`MEM('o046524, 16'o000000);
`MEM('o046526, 16'o000000);
`MEM('o046530, 16'o000000);
`MEM('o046532, 16'o000000);
`MEM('o046534, 16'o000000);
`MEM('o046536, 16'o000000);
`MEM('o046540, 16'o000000);
`MEM('o046542, 16'o000000);
`MEM('o046544, 16'o000000);
`MEM('o046546, 16'o000000);
`MEM('o046550, 16'o000000);
`MEM('o046552, 16'o000000);
`MEM('o046554, 16'o000000);
`MEM('o046556, 16'o000000);
`MEM('o046560, 16'o000000);
`MEM('o046562, 16'o000000);
`MEM('o046564, 16'o000000);
`MEM('o046566, 16'o000000);
`MEM('o046570, 16'o000000);
`MEM('o046572, 16'o000000);
`MEM('o046574, 16'o000000);
`MEM('o046576, 16'o000000);
`MEM('o046600, 16'o000000);
`MEM('o046602, 16'o000000);
`MEM('o046604, 16'o000000);
`MEM('o046606, 16'o000000);
`MEM('o046610, 16'o000000);
`MEM('o046612, 16'o000000);
`MEM('o046614, 16'o000000);
`MEM('o046616, 16'o000000);
`MEM('o046620, 16'o000000);
`MEM('o046622, 16'o000000);
`MEM('o046624, 16'o000000);
`MEM('o046626, 16'o000000);
`MEM('o046630, 16'o000000);
`MEM('o046632, 16'o000000);
`MEM('o046634, 16'o000000);
`MEM('o046636, 16'o000000);
`MEM('o046640, 16'o000000);
`MEM('o046642, 16'o000000);
`MEM('o046644, 16'o000000);
`MEM('o046646, 16'o000000);
`MEM('o046650, 16'o000000);
`MEM('o046652, 16'o000000);
`MEM('o046654, 16'o000000);
`MEM('o046656, 16'o000000);
`MEM('o046660, 16'o000000);
`MEM('o046662, 16'o000000);
`MEM('o046664, 16'o000000);
`MEM('o046666, 16'o000000);
`MEM('o046670, 16'o000000);
`MEM('o046672, 16'o000000);
`MEM('o046674, 16'o000000);
`MEM('o046676, 16'o000000);
`MEM('o046700, 16'o000000);
`MEM('o046702, 16'o000000);
`MEM('o046704, 16'o000000);
`MEM('o046706, 16'o000000);
`MEM('o046710, 16'o000000);
`MEM('o046712, 16'o000000);
`MEM('o046714, 16'o000000);
`MEM('o046716, 16'o000000);
`MEM('o046720, 16'o000000);
`MEM('o046722, 16'o000000);
`MEM('o046724, 16'o000000);
`MEM('o046726, 16'o000000);
`MEM('o046730, 16'o000000);
`MEM('o046732, 16'o000000);
`MEM('o046734, 16'o000000);
`MEM('o046736, 16'o000000);
`MEM('o046740, 16'o000000);
`MEM('o046742, 16'o000000);
`MEM('o046744, 16'o000000);
`MEM('o046746, 16'o000000);
`MEM('o046750, 16'o000000);
`MEM('o046752, 16'o000000);
`MEM('o046754, 16'o000000);
`MEM('o046756, 16'o000000);
`MEM('o046760, 16'o000000);
`MEM('o046762, 16'o000000);
`MEM('o046764, 16'o000000);
`MEM('o046766, 16'o000000);
`MEM('o046770, 16'o000000);
`MEM('o046772, 16'o000000);
`MEM('o046774, 16'o000000);
`MEM('o046776, 16'o000000);
`MEM('o047000, 16'o000000);
`MEM('o047002, 16'o000000);
`MEM('o047004, 16'o000000);
`MEM('o047006, 16'o000000);
`MEM('o047010, 16'o000000);
`MEM('o047012, 16'o000000);
`MEM('o047014, 16'o000000);
`MEM('o047016, 16'o000000);
`MEM('o047020, 16'o000000);
`MEM('o047022, 16'o000000);
`MEM('o047024, 16'o000000);
`MEM('o047026, 16'o000000);
`MEM('o047030, 16'o000000);
`MEM('o047032, 16'o000000);
`MEM('o047034, 16'o000000);
`MEM('o047036, 16'o000000);
`MEM('o047040, 16'o000000);
`MEM('o047042, 16'o000000);
`MEM('o047044, 16'o000000);
`MEM('o047046, 16'o000000);
`MEM('o047050, 16'o000000);
`MEM('o047052, 16'o000000);
`MEM('o047054, 16'o000000);
`MEM('o047056, 16'o000000);
`MEM('o047060, 16'o000000);
`MEM('o047062, 16'o000000);
`MEM('o047064, 16'o000000);
`MEM('o047066, 16'o000000);
`MEM('o047070, 16'o000000);
`MEM('o047072, 16'o000000);
`MEM('o047074, 16'o000000);
`MEM('o047076, 16'o000000);
`MEM('o047100, 16'o000000);
`MEM('o047102, 16'o000000);
`MEM('o047104, 16'o000000);
`MEM('o047106, 16'o000000);
`MEM('o047110, 16'o000000);
`MEM('o047112, 16'o000000);
`MEM('o047114, 16'o000000);
`MEM('o047116, 16'o000000);
`MEM('o047120, 16'o000000);
`MEM('o047122, 16'o000000);
`MEM('o047124, 16'o000000);
`MEM('o047126, 16'o000000);
`MEM('o047130, 16'o000000);
`MEM('o047132, 16'o000000);
`MEM('o047134, 16'o000000);
`MEM('o047136, 16'o000000);
`MEM('o047140, 16'o000000);
`MEM('o047142, 16'o000000);
`MEM('o047144, 16'o000000);
`MEM('o047146, 16'o000000);
`MEM('o047150, 16'o000000);
`MEM('o047152, 16'o000000);
`MEM('o047154, 16'o000000);
`MEM('o047156, 16'o000000);
`MEM('o047160, 16'o000000);
`MEM('o047162, 16'o000000);
`MEM('o047164, 16'o000000);
`MEM('o047166, 16'o000000);
`MEM('o047170, 16'o000000);
`MEM('o047172, 16'o000000);
`MEM('o047174, 16'o000000);
`MEM('o047176, 16'o000000);
`MEM('o047200, 16'o000000);
`MEM('o047202, 16'o000000);
`MEM('o047204, 16'o000000);
`MEM('o047206, 16'o000000);
`MEM('o047210, 16'o000000);
`MEM('o047212, 16'o000000);
`MEM('o047214, 16'o000000);
`MEM('o047216, 16'o000000);
`MEM('o047220, 16'o000000);
`MEM('o047222, 16'o000000);
`MEM('o047224, 16'o000000);
`MEM('o047226, 16'o000000);
`MEM('o047230, 16'o000000);
`MEM('o047232, 16'o000000);
`MEM('o047234, 16'o000000);
`MEM('o047236, 16'o000000);
`MEM('o047240, 16'o000000);
`MEM('o047242, 16'o000000);
`MEM('o047244, 16'o000000);
`MEM('o047246, 16'o000000);
`MEM('o047250, 16'o000000);
`MEM('o047252, 16'o000000);
`MEM('o047254, 16'o000000);
`MEM('o047256, 16'o000000);
`MEM('o047260, 16'o000000);
`MEM('o047262, 16'o000000);
`MEM('o047264, 16'o000000);
`MEM('o047266, 16'o000000);
`MEM('o047270, 16'o000000);
`MEM('o047272, 16'o000000);
`MEM('o047274, 16'o000000);
`MEM('o047276, 16'o000000);
`MEM('o047300, 16'o000000);
`MEM('o047302, 16'o000000);
`MEM('o047304, 16'o000000);
`MEM('o047306, 16'o000000);
`MEM('o047310, 16'o000000);
`MEM('o047312, 16'o000000);
`MEM('o047314, 16'o000000);
`MEM('o047316, 16'o000000);
`MEM('o047320, 16'o000000);
`MEM('o047322, 16'o000000);
`MEM('o047324, 16'o000000);
`MEM('o047326, 16'o000000);
`MEM('o047330, 16'o000000);
`MEM('o047332, 16'o000000);
`MEM('o047334, 16'o000000);
`MEM('o047336, 16'o000000);
`MEM('o047340, 16'o000000);
`MEM('o047342, 16'o000000);
`MEM('o047344, 16'o000000);
`MEM('o047346, 16'o000000);
`MEM('o047350, 16'o000000);
`MEM('o047352, 16'o000000);
`MEM('o047354, 16'o000000);
`MEM('o047356, 16'o000000);
`MEM('o047360, 16'o000000);
`MEM('o047362, 16'o000000);
`MEM('o047364, 16'o000000);
`MEM('o047366, 16'o000000);
`MEM('o047370, 16'o000000);
`MEM('o047372, 16'o000000);
`MEM('o047374, 16'o000000);
`MEM('o047376, 16'o000000);
`MEM('o047400, 16'o000000);
`MEM('o047402, 16'o000000);
`MEM('o047404, 16'o000000);
`MEM('o047406, 16'o000000);
`MEM('o047410, 16'o000000);
`MEM('o047412, 16'o000000);
`MEM('o047414, 16'o000000);
`MEM('o047416, 16'o000000);
`MEM('o047420, 16'o000000);
`MEM('o047422, 16'o000000);
`MEM('o047424, 16'o000000);
`MEM('o047426, 16'o000000);
`MEM('o047430, 16'o000000);
`MEM('o047432, 16'o000000);
`MEM('o047434, 16'o000000);
`MEM('o047436, 16'o000000);
`MEM('o047440, 16'o000000);
`MEM('o047442, 16'o000000);
`MEM('o047444, 16'o000000);
`MEM('o047446, 16'o000000);
`MEM('o047450, 16'o000000);
`MEM('o047452, 16'o000000);
`MEM('o047454, 16'o000000);
`MEM('o047456, 16'o000000);
`MEM('o047460, 16'o000000);
`MEM('o047462, 16'o000000);
`MEM('o047464, 16'o000000);
`MEM('o047466, 16'o000000);
`MEM('o047470, 16'o000000);
`MEM('o047472, 16'o000000);
`MEM('o047474, 16'o000000);
`MEM('o047476, 16'o000000);
`MEM('o047500, 16'o000000);
`MEM('o047502, 16'o000000);
`MEM('o047504, 16'o000000);
`MEM('o047506, 16'o000000);
`MEM('o047510, 16'o000000);
`MEM('o047512, 16'o000000);
`MEM('o047514, 16'o000000);
`MEM('o047516, 16'o000000);
`MEM('o047520, 16'o000000);
`MEM('o047522, 16'o000000);
`MEM('o047524, 16'o000000);
`MEM('o047526, 16'o000000);
`MEM('o047530, 16'o000000);
`MEM('o047532, 16'o000000);
`MEM('o047534, 16'o000000);
`MEM('o047536, 16'o000000);
`MEM('o047540, 16'o000000);
`MEM('o047542, 16'o000000);
`MEM('o047544, 16'o000000);
`MEM('o047546, 16'o000000);
`MEM('o047550, 16'o000000);
`MEM('o047552, 16'o000000);
`MEM('o047554, 16'o000000);
`MEM('o047556, 16'o000000);
`MEM('o047560, 16'o000000);
`MEM('o047562, 16'o000000);
`MEM('o047564, 16'o000000);
`MEM('o047566, 16'o000000);
`MEM('o047570, 16'o000000);
`MEM('o047572, 16'o000000);
`MEM('o047574, 16'o000000);
`MEM('o047576, 16'o000000);
`MEM('o047600, 16'o000000);
`MEM('o047602, 16'o000000);
`MEM('o047604, 16'o000000);
`MEM('o047606, 16'o000000);
`MEM('o047610, 16'o000000);
`MEM('o047612, 16'o000000);
`MEM('o047614, 16'o000000);
`MEM('o047616, 16'o000000);
`MEM('o047620, 16'o000000);
`MEM('o047622, 16'o000000);
`MEM('o047624, 16'o000000);
`MEM('o047626, 16'o000000);
`MEM('o047630, 16'o000000);
`MEM('o047632, 16'o000000);
`MEM('o047634, 16'o000000);
`MEM('o047636, 16'o000000);
`MEM('o047640, 16'o000000);
`MEM('o047642, 16'o000000);
`MEM('o047644, 16'o000000);
`MEM('o047646, 16'o000000);
`MEM('o047650, 16'o000000);
`MEM('o047652, 16'o000000);
`MEM('o047654, 16'o000000);
`MEM('o047656, 16'o000000);
`MEM('o047660, 16'o000000);
`MEM('o047662, 16'o000000);
`MEM('o047664, 16'o000000);
`MEM('o047666, 16'o000000);
`MEM('o047670, 16'o000000);
`MEM('o047672, 16'o000000);
`MEM('o047674, 16'o000000);
`MEM('o047676, 16'o000000);
`MEM('o047700, 16'o000000);
`MEM('o047702, 16'o000000);
`MEM('o047704, 16'o000000);
`MEM('o047706, 16'o000000);
`MEM('o047710, 16'o000000);
`MEM('o047712, 16'o000000);
`MEM('o047714, 16'o000000);
`MEM('o047716, 16'o000000);
`MEM('o047720, 16'o000000);
`MEM('o047722, 16'o000000);
`MEM('o047724, 16'o000000);
`MEM('o047726, 16'o000000);
`MEM('o047730, 16'o000000);
`MEM('o047732, 16'o000000);
`MEM('o047734, 16'o000000);
`MEM('o047736, 16'o000000);
`MEM('o047740, 16'o000000);
`MEM('o047742, 16'o000000);
`MEM('o047744, 16'o000000);
`MEM('o047746, 16'o000000);
`MEM('o047750, 16'o000000);
`MEM('o047752, 16'o000000);
`MEM('o047754, 16'o000000);
`MEM('o047756, 16'o000000);
`MEM('o047760, 16'o000000);
`MEM('o047762, 16'o000000);
`MEM('o047764, 16'o000000);
`MEM('o047766, 16'o000000);
`MEM('o047770, 16'o000000);
`MEM('o047772, 16'o000000);
`MEM('o047774, 16'o000000);
`MEM('o047776, 16'o000000);
`MEM('o050000, 16'o000000);
`MEM('o050002, 16'o000000);
`MEM('o050004, 16'o000000);
`MEM('o050006, 16'o000000);
`MEM('o050010, 16'o000000);
`MEM('o050012, 16'o000000);
`MEM('o050014, 16'o000000);
`MEM('o050016, 16'o000000);
`MEM('o050020, 16'o000000);
`MEM('o050022, 16'o000000);
`MEM('o050024, 16'o000000);
`MEM('o050026, 16'o000000);
`MEM('o050030, 16'o000000);
`MEM('o050032, 16'o000000);
`MEM('o050034, 16'o000000);
`MEM('o050036, 16'o000000);
`MEM('o050040, 16'o000000);
`MEM('o050042, 16'o000000);
`MEM('o050044, 16'o000000);
`MEM('o050046, 16'o000000);
`MEM('o050050, 16'o000000);
`MEM('o050052, 16'o000000);
`MEM('o050054, 16'o000000);
`MEM('o050056, 16'o000000);
`MEM('o050060, 16'o000000);
`MEM('o050062, 16'o000000);
`MEM('o050064, 16'o000000);
`MEM('o050066, 16'o000000);
`MEM('o050070, 16'o000000);
`MEM('o050072, 16'o000000);
`MEM('o050074, 16'o000000);
`MEM('o050076, 16'o000000);
`MEM('o050100, 16'o000000);
`MEM('o050102, 16'o000000);
`MEM('o050104, 16'o000000);
`MEM('o050106, 16'o000000);
`MEM('o050110, 16'o000000);
`MEM('o050112, 16'o000000);
`MEM('o050114, 16'o000000);
`MEM('o050116, 16'o000000);
`MEM('o050120, 16'o000000);
`MEM('o050122, 16'o000000);
`MEM('o050124, 16'o000000);
`MEM('o050126, 16'o000000);
`MEM('o050130, 16'o000000);
`MEM('o050132, 16'o000000);
`MEM('o050134, 16'o000000);
`MEM('o050136, 16'o000000);
`MEM('o050140, 16'o000000);
`MEM('o050142, 16'o000000);
`MEM('o050144, 16'o000000);
`MEM('o050146, 16'o000000);
`MEM('o050150, 16'o000000);
`MEM('o050152, 16'o000000);
`MEM('o050154, 16'o000000);
`MEM('o050156, 16'o000000);
`MEM('o050160, 16'o000000);
`MEM('o050162, 16'o000000);
`MEM('o050164, 16'o000000);
`MEM('o050166, 16'o000000);
`MEM('o050170, 16'o000000);
`MEM('o050172, 16'o000000);
`MEM('o050174, 16'o000000);
`MEM('o050176, 16'o000000);
`MEM('o050200, 16'o000000);
`MEM('o050202, 16'o000000);
`MEM('o050204, 16'o000000);
`MEM('o050206, 16'o000000);
`MEM('o050210, 16'o000000);
`MEM('o050212, 16'o000000);
`MEM('o050214, 16'o000000);
`MEM('o050216, 16'o000000);
`MEM('o050220, 16'o000000);
`MEM('o050222, 16'o000000);
`MEM('o050224, 16'o000000);
`MEM('o050226, 16'o000000);
`MEM('o050230, 16'o000000);
`MEM('o050232, 16'o000000);
`MEM('o050234, 16'o000000);
`MEM('o050236, 16'o000000);
`MEM('o050240, 16'o000000);
`MEM('o050242, 16'o000000);
`MEM('o050244, 16'o000000);
`MEM('o050246, 16'o000000);
`MEM('o050250, 16'o000000);
`MEM('o050252, 16'o000000);
`MEM('o050254, 16'o000000);
`MEM('o050256, 16'o000000);
`MEM('o050260, 16'o000000);
`MEM('o050262, 16'o000000);
`MEM('o050264, 16'o000000);
`MEM('o050266, 16'o000000);
`MEM('o050270, 16'o000000);
`MEM('o050272, 16'o000000);
`MEM('o050274, 16'o000000);
`MEM('o050276, 16'o000000);
`MEM('o050300, 16'o000000);
`MEM('o050302, 16'o000000);
`MEM('o050304, 16'o000000);
`MEM('o050306, 16'o000000);
`MEM('o050310, 16'o000000);
`MEM('o050312, 16'o000000);
`MEM('o050314, 16'o000000);
`MEM('o050316, 16'o000000);
`MEM('o050320, 16'o000000);
`MEM('o050322, 16'o000000);
`MEM('o050324, 16'o000000);
`MEM('o050326, 16'o000000);
`MEM('o050330, 16'o000000);
`MEM('o050332, 16'o000000);
`MEM('o050334, 16'o000000);
`MEM('o050336, 16'o000000);
`MEM('o050340, 16'o000000);
`MEM('o050342, 16'o000000);
`MEM('o050344, 16'o000000);
`MEM('o050346, 16'o000000);
`MEM('o050350, 16'o000000);
`MEM('o050352, 16'o000000);
`MEM('o050354, 16'o000000);
`MEM('o050356, 16'o000000);
`MEM('o050360, 16'o000000);
`MEM('o050362, 16'o000000);
`MEM('o050364, 16'o000000);
`MEM('o050366, 16'o000000);
`MEM('o050370, 16'o000000);
`MEM('o050372, 16'o000000);
`MEM('o050374, 16'o000000);
`MEM('o050376, 16'o000000);
`MEM('o050400, 16'o000000);
`MEM('o050402, 16'o000000);
`MEM('o050404, 16'o000000);
`MEM('o050406, 16'o000000);
`MEM('o050410, 16'o000000);
`MEM('o050412, 16'o000000);
`MEM('o050414, 16'o000000);
`MEM('o050416, 16'o000000);
`MEM('o050420, 16'o000000);
`MEM('o050422, 16'o000000);
`MEM('o050424, 16'o000000);
`MEM('o050426, 16'o000000);
`MEM('o050430, 16'o000000);
`MEM('o050432, 16'o000000);
`MEM('o050434, 16'o000000);
`MEM('o050436, 16'o000000);
`MEM('o050440, 16'o000000);
`MEM('o050442, 16'o000000);
`MEM('o050444, 16'o000000);
`MEM('o050446, 16'o000000);
`MEM('o050450, 16'o000000);
`MEM('o050452, 16'o000000);
`MEM('o050454, 16'o000000);
`MEM('o050456, 16'o000000);
`MEM('o050460, 16'o000000);
`MEM('o050462, 16'o000000);
`MEM('o050464, 16'o000000);
`MEM('o050466, 16'o000000);
`MEM('o050470, 16'o000000);
`MEM('o050472, 16'o000000);
`MEM('o050474, 16'o000000);
`MEM('o050476, 16'o000000);
`MEM('o050500, 16'o000000);
`MEM('o050502, 16'o000000);
`MEM('o050504, 16'o000000);
`MEM('o050506, 16'o000000);
`MEM('o050510, 16'o000000);
`MEM('o050512, 16'o000000);
`MEM('o050514, 16'o000000);
`MEM('o050516, 16'o000000);
`MEM('o050520, 16'o000000);
`MEM('o050522, 16'o000000);
`MEM('o050524, 16'o000000);
`MEM('o050526, 16'o000000);
`MEM('o050530, 16'o000000);
`MEM('o050532, 16'o000000);
`MEM('o050534, 16'o000000);
`MEM('o050536, 16'o000000);
`MEM('o050540, 16'o000000);
`MEM('o050542, 16'o000000);
`MEM('o050544, 16'o000000);
`MEM('o050546, 16'o000000);
`MEM('o050550, 16'o000000);
`MEM('o050552, 16'o000000);
`MEM('o050554, 16'o000000);
`MEM('o050556, 16'o000000);
`MEM('o050560, 16'o000000);
`MEM('o050562, 16'o000000);
`MEM('o050564, 16'o000000);
`MEM('o050566, 16'o000000);
`MEM('o050570, 16'o000000);
`MEM('o050572, 16'o000000);
`MEM('o050574, 16'o000000);
`MEM('o050576, 16'o000000);
`MEM('o050600, 16'o000000);
`MEM('o050602, 16'o000000);
`MEM('o050604, 16'o000000);
`MEM('o050606, 16'o000000);
`MEM('o050610, 16'o000000);
`MEM('o050612, 16'o000000);
`MEM('o050614, 16'o000000);
`MEM('o050616, 16'o000000);
`MEM('o050620, 16'o000000);
`MEM('o050622, 16'o000000);
`MEM('o050624, 16'o000000);
`MEM('o050626, 16'o000000);
`MEM('o050630, 16'o000000);
`MEM('o050632, 16'o000000);
`MEM('o050634, 16'o000000);
`MEM('o050636, 16'o000000);
`MEM('o050640, 16'o000000);
`MEM('o050642, 16'o000000);
`MEM('o050644, 16'o000000);
`MEM('o050646, 16'o000000);
`MEM('o050650, 16'o000000);
`MEM('o050652, 16'o000000);
`MEM('o050654, 16'o000000);
`MEM('o050656, 16'o000000);
`MEM('o050660, 16'o000000);
`MEM('o050662, 16'o000000);
`MEM('o050664, 16'o000000);
`MEM('o050666, 16'o000000);
`MEM('o050670, 16'o000000);
`MEM('o050672, 16'o000000);
`MEM('o050674, 16'o000000);
`MEM('o050676, 16'o000000);
`MEM('o050700, 16'o000000);
`MEM('o050702, 16'o000000);
`MEM('o050704, 16'o000000);
`MEM('o050706, 16'o000000);
`MEM('o050710, 16'o000000);
`MEM('o050712, 16'o000000);
`MEM('o050714, 16'o000000);
`MEM('o050716, 16'o000000);
`MEM('o050720, 16'o000000);
`MEM('o050722, 16'o000000);
`MEM('o050724, 16'o000000);
`MEM('o050726, 16'o000000);
`MEM('o050730, 16'o000000);
`MEM('o050732, 16'o000000);
`MEM('o050734, 16'o000000);
`MEM('o050736, 16'o000000);
`MEM('o050740, 16'o000000);
`MEM('o050742, 16'o000000);
`MEM('o050744, 16'o000000);
`MEM('o050746, 16'o000000);
`MEM('o050750, 16'o000000);
`MEM('o050752, 16'o000000);
`MEM('o050754, 16'o000000);
`MEM('o050756, 16'o000000);
`MEM('o050760, 16'o000000);
`MEM('o050762, 16'o000000);
`MEM('o050764, 16'o000000);
`MEM('o050766, 16'o000000);
`MEM('o050770, 16'o000000);
`MEM('o050772, 16'o000000);
`MEM('o050774, 16'o000000);
`MEM('o050776, 16'o000000);
`MEM('o051000, 16'o000000);
`MEM('o051002, 16'o000000);
`MEM('o051004, 16'o000000);
`MEM('o051006, 16'o000000);
`MEM('o051010, 16'o000000);
`MEM('o051012, 16'o000000);
`MEM('o051014, 16'o000000);
`MEM('o051016, 16'o000000);
`MEM('o051020, 16'o000000);
`MEM('o051022, 16'o000000);
`MEM('o051024, 16'o000000);
`MEM('o051026, 16'o000000);
`MEM('o051030, 16'o000000);
`MEM('o051032, 16'o000000);
`MEM('o051034, 16'o000000);
`MEM('o051036, 16'o000000);
`MEM('o051040, 16'o000000);
`MEM('o051042, 16'o000000);
`MEM('o051044, 16'o000000);
`MEM('o051046, 16'o000000);
`MEM('o051050, 16'o000000);
`MEM('o051052, 16'o000000);
`MEM('o051054, 16'o000000);
`MEM('o051056, 16'o000000);
`MEM('o051060, 16'o000000);
`MEM('o051062, 16'o000000);
`MEM('o051064, 16'o000000);
`MEM('o051066, 16'o000000);
`MEM('o051070, 16'o000000);
`MEM('o051072, 16'o000000);
`MEM('o051074, 16'o000000);
`MEM('o051076, 16'o000000);
`MEM('o051100, 16'o000000);
`MEM('o051102, 16'o000000);
`MEM('o051104, 16'o000000);
`MEM('o051106, 16'o000000);
`MEM('o051110, 16'o000000);
`MEM('o051112, 16'o000000);
`MEM('o051114, 16'o000000);
`MEM('o051116, 16'o000000);
`MEM('o051120, 16'o000000);
`MEM('o051122, 16'o000000);
`MEM('o051124, 16'o000000);
`MEM('o051126, 16'o000000);
`MEM('o051130, 16'o000000);
`MEM('o051132, 16'o000000);
`MEM('o051134, 16'o000000);
`MEM('o051136, 16'o000000);
`MEM('o051140, 16'o000000);
`MEM('o051142, 16'o000000);
`MEM('o051144, 16'o000000);
`MEM('o051146, 16'o000000);
`MEM('o051150, 16'o000000);
`MEM('o051152, 16'o000000);
`MEM('o051154, 16'o000000);
`MEM('o051156, 16'o000000);
`MEM('o051160, 16'o000000);
`MEM('o051162, 16'o000000);
`MEM('o051164, 16'o000000);
`MEM('o051166, 16'o000000);
`MEM('o051170, 16'o000000);
`MEM('o051172, 16'o000000);
`MEM('o051174, 16'o000000);
`MEM('o051176, 16'o000000);
`MEM('o051200, 16'o000000);
`MEM('o051202, 16'o000000);
`MEM('o051204, 16'o000000);
`MEM('o051206, 16'o000000);
`MEM('o051210, 16'o000000);
`MEM('o051212, 16'o000000);
`MEM('o051214, 16'o000000);
`MEM('o051216, 16'o000000);
`MEM('o051220, 16'o000000);
`MEM('o051222, 16'o000000);
`MEM('o051224, 16'o000000);
`MEM('o051226, 16'o000000);
`MEM('o051230, 16'o000000);
`MEM('o051232, 16'o000000);
`MEM('o051234, 16'o000000);
`MEM('o051236, 16'o000000);
`MEM('o051240, 16'o000000);
`MEM('o051242, 16'o000000);
`MEM('o051244, 16'o000000);
`MEM('o051246, 16'o000000);
`MEM('o051250, 16'o000000);
`MEM('o051252, 16'o000000);
`MEM('o051254, 16'o000000);
`MEM('o051256, 16'o000000);
`MEM('o051260, 16'o000000);
`MEM('o051262, 16'o000000);
`MEM('o051264, 16'o000000);
`MEM('o051266, 16'o000000);
`MEM('o051270, 16'o000000);
`MEM('o051272, 16'o000000);
`MEM('o051274, 16'o000000);
`MEM('o051276, 16'o000000);
`MEM('o051300, 16'o000000);
`MEM('o051302, 16'o000000);
`MEM('o051304, 16'o000000);
`MEM('o051306, 16'o000000);
`MEM('o051310, 16'o000000);
`MEM('o051312, 16'o000000);
`MEM('o051314, 16'o000000);
`MEM('o051316, 16'o000000);
`MEM('o051320, 16'o000000);
`MEM('o051322, 16'o000000);
`MEM('o051324, 16'o000000);
`MEM('o051326, 16'o000000);
`MEM('o051330, 16'o000000);
`MEM('o051332, 16'o000000);
`MEM('o051334, 16'o000000);
`MEM('o051336, 16'o000000);
`MEM('o051340, 16'o000000);
`MEM('o051342, 16'o000000);
`MEM('o051344, 16'o000000);
`MEM('o051346, 16'o000000);
`MEM('o051350, 16'o000000);
`MEM('o051352, 16'o000000);
`MEM('o051354, 16'o000000);
`MEM('o051356, 16'o000000);
`MEM('o051360, 16'o000000);
`MEM('o051362, 16'o000000);
`MEM('o051364, 16'o000000);
`MEM('o051366, 16'o000000);
`MEM('o051370, 16'o000000);
`MEM('o051372, 16'o000000);
`MEM('o051374, 16'o000000);
`MEM('o051376, 16'o000000);
`MEM('o051400, 16'o000000);
`MEM('o051402, 16'o000000);
`MEM('o051404, 16'o000000);
`MEM('o051406, 16'o000000);
`MEM('o051410, 16'o000000);
`MEM('o051412, 16'o000000);
`MEM('o051414, 16'o000000);
`MEM('o051416, 16'o000000);
`MEM('o051420, 16'o000000);
`MEM('o051422, 16'o000000);
`MEM('o051424, 16'o000000);
`MEM('o051426, 16'o000000);
`MEM('o051430, 16'o000000);
`MEM('o051432, 16'o000000);
`MEM('o051434, 16'o000000);
`MEM('o051436, 16'o000000);
`MEM('o051440, 16'o000000);
`MEM('o051442, 16'o000000);
`MEM('o051444, 16'o000000);
`MEM('o051446, 16'o000000);
`MEM('o051450, 16'o000000);
`MEM('o051452, 16'o000000);
`MEM('o051454, 16'o000000);
`MEM('o051456, 16'o000000);
`MEM('o051460, 16'o000000);
`MEM('o051462, 16'o000000);
`MEM('o051464, 16'o000000);
`MEM('o051466, 16'o000000);
`MEM('o051470, 16'o000000);
`MEM('o051472, 16'o000000);
`MEM('o051474, 16'o000000);
`MEM('o051476, 16'o000000);
`MEM('o051500, 16'o000000);
`MEM('o051502, 16'o000000);
`MEM('o051504, 16'o000000);
`MEM('o051506, 16'o000000);
`MEM('o051510, 16'o000000);
`MEM('o051512, 16'o000000);
`MEM('o051514, 16'o000000);
`MEM('o051516, 16'o000000);
`MEM('o051520, 16'o000000);
`MEM('o051522, 16'o000000);
`MEM('o051524, 16'o000000);
`MEM('o051526, 16'o000000);
`MEM('o051530, 16'o000000);
`MEM('o051532, 16'o000000);
`MEM('o051534, 16'o000000);
`MEM('o051536, 16'o000000);
`MEM('o051540, 16'o000000);
`MEM('o051542, 16'o000000);
`MEM('o051544, 16'o000000);
`MEM('o051546, 16'o000000);
`MEM('o051550, 16'o000000);
`MEM('o051552, 16'o000000);
`MEM('o051554, 16'o000000);
`MEM('o051556, 16'o000000);
`MEM('o051560, 16'o000000);
`MEM('o051562, 16'o000000);
`MEM('o051564, 16'o000000);
`MEM('o051566, 16'o000000);
`MEM('o051570, 16'o000000);
`MEM('o051572, 16'o000000);
`MEM('o051574, 16'o000000);
`MEM('o051576, 16'o000000);
`MEM('o051600, 16'o000000);
`MEM('o051602, 16'o000000);
`MEM('o051604, 16'o000000);
`MEM('o051606, 16'o000000);
`MEM('o051610, 16'o000000);
`MEM('o051612, 16'o000000);
`MEM('o051614, 16'o000000);
`MEM('o051616, 16'o000000);
`MEM('o051620, 16'o000000);
`MEM('o051622, 16'o000000);
`MEM('o051624, 16'o000000);
`MEM('o051626, 16'o000000);
`MEM('o051630, 16'o000000);
`MEM('o051632, 16'o000000);
`MEM('o051634, 16'o000000);
`MEM('o051636, 16'o000000);
`MEM('o051640, 16'o000000);
`MEM('o051642, 16'o000000);
`MEM('o051644, 16'o000000);
`MEM('o051646, 16'o000000);
`MEM('o051650, 16'o000000);
`MEM('o051652, 16'o000000);
`MEM('o051654, 16'o000000);
`MEM('o051656, 16'o000000);
`MEM('o051660, 16'o000000);
`MEM('o051662, 16'o000000);
`MEM('o051664, 16'o000000);
`MEM('o051666, 16'o000000);
`MEM('o051670, 16'o000000);
`MEM('o051672, 16'o000000);
`MEM('o051674, 16'o000000);
`MEM('o051676, 16'o000000);
`MEM('o051700, 16'o000000);
`MEM('o051702, 16'o000000);
`MEM('o051704, 16'o000000);
`MEM('o051706, 16'o000000);
`MEM('o051710, 16'o000000);
`MEM('o051712, 16'o000000);
`MEM('o051714, 16'o000000);
`MEM('o051716, 16'o000000);
`MEM('o051720, 16'o000000);
`MEM('o051722, 16'o000000);
`MEM('o051724, 16'o000000);
`MEM('o051726, 16'o000000);
`MEM('o051730, 16'o000000);
`MEM('o051732, 16'o000000);
`MEM('o051734, 16'o000000);
`MEM('o051736, 16'o000000);
`MEM('o051740, 16'o000000);
`MEM('o051742, 16'o000000);
`MEM('o051744, 16'o000000);
`MEM('o051746, 16'o000000);
`MEM('o051750, 16'o000000);
`MEM('o051752, 16'o000000);
`MEM('o051754, 16'o000000);
`MEM('o051756, 16'o000000);
`MEM('o051760, 16'o000000);
`MEM('o051762, 16'o000000);
`MEM('o051764, 16'o000000);
`MEM('o051766, 16'o000000);
`MEM('o051770, 16'o000000);
`MEM('o051772, 16'o000000);
`MEM('o051774, 16'o000000);
`MEM('o051776, 16'o000000);
`MEM('o052000, 16'o000000);
`MEM('o052002, 16'o000000);
`MEM('o052004, 16'o000000);
`MEM('o052006, 16'o000000);
`MEM('o052010, 16'o000000);
`MEM('o052012, 16'o000000);
`MEM('o052014, 16'o000000);
`MEM('o052016, 16'o000000);
`MEM('o052020, 16'o000000);
`MEM('o052022, 16'o000000);
`MEM('o052024, 16'o000000);
`MEM('o052026, 16'o000000);
`MEM('o052030, 16'o000000);
`MEM('o052032, 16'o000000);
`MEM('o052034, 16'o000000);
`MEM('o052036, 16'o000000);
`MEM('o052040, 16'o000000);
`MEM('o052042, 16'o000000);
`MEM('o052044, 16'o000000);
`MEM('o052046, 16'o000000);
`MEM('o052050, 16'o000000);
`MEM('o052052, 16'o000000);
`MEM('o052054, 16'o000000);
`MEM('o052056, 16'o000000);
`MEM('o052060, 16'o000000);
`MEM('o052062, 16'o000000);
`MEM('o052064, 16'o000000);
`MEM('o052066, 16'o000000);
`MEM('o052070, 16'o000000);
`MEM('o052072, 16'o000000);
`MEM('o052074, 16'o000000);
`MEM('o052076, 16'o000000);
`MEM('o052100, 16'o000000);
`MEM('o052102, 16'o000000);
`MEM('o052104, 16'o000000);
`MEM('o052106, 16'o000000);
`MEM('o052110, 16'o000000);
`MEM('o052112, 16'o000000);
`MEM('o052114, 16'o000000);
`MEM('o052116, 16'o000000);
`MEM('o052120, 16'o000000);
`MEM('o052122, 16'o000000);
`MEM('o052124, 16'o000000);
`MEM('o052126, 16'o000000);
`MEM('o052130, 16'o000000);
`MEM('o052132, 16'o000000);
`MEM('o052134, 16'o000000);
`MEM('o052136, 16'o000000);
`MEM('o052140, 16'o000000);
`MEM('o052142, 16'o000000);
`MEM('o052144, 16'o000000);
`MEM('o052146, 16'o000000);
`MEM('o052150, 16'o000000);
`MEM('o052152, 16'o000000);
`MEM('o052154, 16'o000000);
`MEM('o052156, 16'o000000);
`MEM('o052160, 16'o000000);
`MEM('o052162, 16'o000000);
`MEM('o052164, 16'o000000);
`MEM('o052166, 16'o000000);
`MEM('o052170, 16'o000000);
`MEM('o052172, 16'o000000);
`MEM('o052174, 16'o000000);
`MEM('o052176, 16'o000000);
`MEM('o052200, 16'o000000);
`MEM('o052202, 16'o000000);
`MEM('o052204, 16'o000000);
`MEM('o052206, 16'o000000);
`MEM('o052210, 16'o000000);
`MEM('o052212, 16'o000000);
`MEM('o052214, 16'o000000);
`MEM('o052216, 16'o000000);
`MEM('o052220, 16'o000000);
`MEM('o052222, 16'o000000);
`MEM('o052224, 16'o000000);
`MEM('o052226, 16'o000000);
`MEM('o052230, 16'o000000);
`MEM('o052232, 16'o000000);
`MEM('o052234, 16'o000000);
`MEM('o052236, 16'o000000);
`MEM('o052240, 16'o000000);
`MEM('o052242, 16'o000000);
`MEM('o052244, 16'o000000);
`MEM('o052246, 16'o000000);
`MEM('o052250, 16'o000000);
`MEM('o052252, 16'o000000);
`MEM('o052254, 16'o000000);
`MEM('o052256, 16'o000000);
`MEM('o052260, 16'o000000);
`MEM('o052262, 16'o000000);
`MEM('o052264, 16'o000000);
`MEM('o052266, 16'o000000);
`MEM('o052270, 16'o000000);
`MEM('o052272, 16'o000000);
`MEM('o052274, 16'o000000);
`MEM('o052276, 16'o000000);
`MEM('o052300, 16'o000000);
`MEM('o052302, 16'o000000);
`MEM('o052304, 16'o000000);
`MEM('o052306, 16'o000000);
`MEM('o052310, 16'o000000);
`MEM('o052312, 16'o000000);
`MEM('o052314, 16'o000000);
`MEM('o052316, 16'o000000);
`MEM('o052320, 16'o000000);
`MEM('o052322, 16'o000000);
`MEM('o052324, 16'o000000);
`MEM('o052326, 16'o000000);
`MEM('o052330, 16'o000000);
`MEM('o052332, 16'o000000);
`MEM('o052334, 16'o000000);
`MEM('o052336, 16'o000000);
`MEM('o052340, 16'o000000);
`MEM('o052342, 16'o000000);
`MEM('o052344, 16'o000000);
`MEM('o052346, 16'o000000);
`MEM('o052350, 16'o000000);
`MEM('o052352, 16'o000000);
`MEM('o052354, 16'o000000);
`MEM('o052356, 16'o000000);
`MEM('o052360, 16'o000000);
`MEM('o052362, 16'o000000);
`MEM('o052364, 16'o000000);
`MEM('o052366, 16'o000000);
`MEM('o052370, 16'o000000);
`MEM('o052372, 16'o000000);
`MEM('o052374, 16'o000000);
`MEM('o052376, 16'o000000);
`MEM('o052400, 16'o000000);
`MEM('o052402, 16'o000000);
`MEM('o052404, 16'o000000);
`MEM('o052406, 16'o000000);
`MEM('o052410, 16'o000000);
`MEM('o052412, 16'o000000);
`MEM('o052414, 16'o000000);
`MEM('o052416, 16'o000000);
`MEM('o052420, 16'o000000);
`MEM('o052422, 16'o000000);
`MEM('o052424, 16'o000000);
`MEM('o052426, 16'o000000);
`MEM('o052430, 16'o000000);
`MEM('o052432, 16'o000000);
`MEM('o052434, 16'o000000);
`MEM('o052436, 16'o000000);
`MEM('o052440, 16'o000000);
`MEM('o052442, 16'o000000);
`MEM('o052444, 16'o000000);
`MEM('o052446, 16'o000000);
`MEM('o052450, 16'o000000);
`MEM('o052452, 16'o000000);
`MEM('o052454, 16'o000000);
`MEM('o052456, 16'o000000);
`MEM('o052460, 16'o000000);
`MEM('o052462, 16'o000000);
`MEM('o052464, 16'o000000);
`MEM('o052466, 16'o000000);
`MEM('o052470, 16'o000000);
`MEM('o052472, 16'o000000);
`MEM('o052474, 16'o000000);
`MEM('o052476, 16'o000000);
`MEM('o052500, 16'o000000);
`MEM('o052502, 16'o000000);
`MEM('o052504, 16'o000000);
`MEM('o052506, 16'o000000);
`MEM('o052510, 16'o000000);
`MEM('o052512, 16'o000000);
`MEM('o052514, 16'o000000);
`MEM('o052516, 16'o000000);
`MEM('o052520, 16'o000000);
`MEM('o052522, 16'o000000);
`MEM('o052524, 16'o000000);
`MEM('o052526, 16'o000000);
`MEM('o052530, 16'o000000);
`MEM('o052532, 16'o000000);
`MEM('o052534, 16'o000000);
`MEM('o052536, 16'o000000);
`MEM('o052540, 16'o000000);
`MEM('o052542, 16'o000000);
`MEM('o052544, 16'o000000);
`MEM('o052546, 16'o000000);
`MEM('o052550, 16'o000000);
`MEM('o052552, 16'o000000);
`MEM('o052554, 16'o000000);
`MEM('o052556, 16'o000000);
`MEM('o052560, 16'o000000);
`MEM('o052562, 16'o000000);
`MEM('o052564, 16'o000000);
`MEM('o052566, 16'o000000);
`MEM('o052570, 16'o000000);
`MEM('o052572, 16'o000000);
`MEM('o052574, 16'o000000);
`MEM('o052576, 16'o000000);
`MEM('o052600, 16'o000000);
`MEM('o052602, 16'o000000);
`MEM('o052604, 16'o000000);
`MEM('o052606, 16'o000000);
`MEM('o052610, 16'o000000);
`MEM('o052612, 16'o000000);
`MEM('o052614, 16'o000000);
`MEM('o052616, 16'o000000);
`MEM('o052620, 16'o000000);
`MEM('o052622, 16'o000000);
`MEM('o052624, 16'o000000);
`MEM('o052626, 16'o000000);
`MEM('o052630, 16'o000000);
`MEM('o052632, 16'o000000);
`MEM('o052634, 16'o000000);
`MEM('o052636, 16'o000000);
`MEM('o052640, 16'o000000);
`MEM('o052642, 16'o000000);
`MEM('o052644, 16'o000000);
`MEM('o052646, 16'o000000);
`MEM('o052650, 16'o000000);
`MEM('o052652, 16'o000000);
`MEM('o052654, 16'o000000);
`MEM('o052656, 16'o000000);
`MEM('o052660, 16'o000000);
`MEM('o052662, 16'o000000);
`MEM('o052664, 16'o000000);
`MEM('o052666, 16'o000000);
`MEM('o052670, 16'o000000);
`MEM('o052672, 16'o000000);
`MEM('o052674, 16'o000000);
`MEM('o052676, 16'o000000);
`MEM('o052700, 16'o000000);
`MEM('o052702, 16'o000000);
`MEM('o052704, 16'o000000);
`MEM('o052706, 16'o000000);
`MEM('o052710, 16'o000000);
`MEM('o052712, 16'o000000);
`MEM('o052714, 16'o000000);
`MEM('o052716, 16'o000000);
`MEM('o052720, 16'o000000);
`MEM('o052722, 16'o000000);
`MEM('o052724, 16'o000000);
`MEM('o052726, 16'o000000);
`MEM('o052730, 16'o000000);
`MEM('o052732, 16'o000000);
`MEM('o052734, 16'o000000);
`MEM('o052736, 16'o000000);
`MEM('o052740, 16'o000000);
`MEM('o052742, 16'o000000);
`MEM('o052744, 16'o000000);
`MEM('o052746, 16'o000000);
`MEM('o052750, 16'o000000);
`MEM('o052752, 16'o000000);
`MEM('o052754, 16'o000000);
`MEM('o052756, 16'o000000);
`MEM('o052760, 16'o000000);
`MEM('o052762, 16'o000000);
`MEM('o052764, 16'o000000);
`MEM('o052766, 16'o000000);
`MEM('o052770, 16'o000000);
`MEM('o052772, 16'o000000);
`MEM('o052774, 16'o000000);
`MEM('o052776, 16'o000000);
`MEM('o053000, 16'o000000);
`MEM('o053002, 16'o000000);
`MEM('o053004, 16'o000000);
`MEM('o053006, 16'o000000);
`MEM('o053010, 16'o000000);
`MEM('o053012, 16'o000000);
`MEM('o053014, 16'o000000);
`MEM('o053016, 16'o000000);
`MEM('o053020, 16'o000000);
`MEM('o053022, 16'o000000);
`MEM('o053024, 16'o000000);
`MEM('o053026, 16'o000000);
`MEM('o053030, 16'o000000);
`MEM('o053032, 16'o000000);
`MEM('o053034, 16'o000000);
`MEM('o053036, 16'o000000);
`MEM('o053040, 16'o000000);
`MEM('o053042, 16'o000000);
`MEM('o053044, 16'o000000);
`MEM('o053046, 16'o000000);
`MEM('o053050, 16'o000000);
`MEM('o053052, 16'o000000);
`MEM('o053054, 16'o000000);
`MEM('o053056, 16'o000000);
`MEM('o053060, 16'o000000);
`MEM('o053062, 16'o000000);
`MEM('o053064, 16'o000000);
`MEM('o053066, 16'o000000);
`MEM('o053070, 16'o000000);
`MEM('o053072, 16'o000000);
`MEM('o053074, 16'o000000);
`MEM('o053076, 16'o000000);
`MEM('o053100, 16'o000000);
`MEM('o053102, 16'o000000);
`MEM('o053104, 16'o000000);
`MEM('o053106, 16'o000000);
`MEM('o053110, 16'o000000);
`MEM('o053112, 16'o000000);
`MEM('o053114, 16'o000000);
`MEM('o053116, 16'o000000);
`MEM('o053120, 16'o000000);
`MEM('o053122, 16'o000000);
`MEM('o053124, 16'o000000);
`MEM('o053126, 16'o000000);
`MEM('o053130, 16'o000000);
`MEM('o053132, 16'o000000);
`MEM('o053134, 16'o000000);
`MEM('o053136, 16'o000000);
`MEM('o053140, 16'o000000);
`MEM('o053142, 16'o000000);
`MEM('o053144, 16'o000000);
`MEM('o053146, 16'o000000);
`MEM('o053150, 16'o000000);
`MEM('o053152, 16'o000000);
`MEM('o053154, 16'o000000);
`MEM('o053156, 16'o000000);
`MEM('o053160, 16'o000000);
`MEM('o053162, 16'o000000);
`MEM('o053164, 16'o000000);
`MEM('o053166, 16'o000000);
`MEM('o053170, 16'o000000);
`MEM('o053172, 16'o000000);
`MEM('o053174, 16'o000000);
`MEM('o053176, 16'o000000);
`MEM('o053200, 16'o000000);
`MEM('o053202, 16'o000000);
`MEM('o053204, 16'o000000);
`MEM('o053206, 16'o000000);
`MEM('o053210, 16'o000000);
`MEM('o053212, 16'o000000);
`MEM('o053214, 16'o000000);
`MEM('o053216, 16'o000000);
`MEM('o053220, 16'o000000);
`MEM('o053222, 16'o000000);
`MEM('o053224, 16'o000000);
`MEM('o053226, 16'o000000);
`MEM('o053230, 16'o000000);
`MEM('o053232, 16'o000000);
`MEM('o053234, 16'o000000);
`MEM('o053236, 16'o000000);
`MEM('o053240, 16'o000000);
`MEM('o053242, 16'o000000);
`MEM('o053244, 16'o000000);
`MEM('o053246, 16'o000000);
`MEM('o053250, 16'o000000);
`MEM('o053252, 16'o000000);
`MEM('o053254, 16'o000000);
`MEM('o053256, 16'o000000);
`MEM('o053260, 16'o000000);
`MEM('o053262, 16'o000000);
`MEM('o053264, 16'o000000);
`MEM('o053266, 16'o000000);
`MEM('o053270, 16'o000000);
`MEM('o053272, 16'o000000);
`MEM('o053274, 16'o000000);
`MEM('o053276, 16'o000000);
`MEM('o053300, 16'o000000);
`MEM('o053302, 16'o000000);
`MEM('o053304, 16'o000000);
`MEM('o053306, 16'o000000);
`MEM('o053310, 16'o000000);
`MEM('o053312, 16'o000000);
`MEM('o053314, 16'o000000);
`MEM('o053316, 16'o000000);
`MEM('o053320, 16'o000000);
`MEM('o053322, 16'o000000);
`MEM('o053324, 16'o000000);
`MEM('o053326, 16'o000000);
`MEM('o053330, 16'o000000);
`MEM('o053332, 16'o000000);
`MEM('o053334, 16'o000000);
`MEM('o053336, 16'o000000);
`MEM('o053340, 16'o000000);
`MEM('o053342, 16'o000000);
`MEM('o053344, 16'o000000);
`MEM('o053346, 16'o000000);
`MEM('o053350, 16'o000000);
`MEM('o053352, 16'o000000);
`MEM('o053354, 16'o000000);
`MEM('o053356, 16'o000000);
`MEM('o053360, 16'o000000);
`MEM('o053362, 16'o000000);
`MEM('o053364, 16'o000000);
`MEM('o053366, 16'o000000);
`MEM('o053370, 16'o000000);
`MEM('o053372, 16'o000000);
`MEM('o053374, 16'o000000);
`MEM('o053376, 16'o000000);
`MEM('o053400, 16'o000000);
`MEM('o053402, 16'o000000);
`MEM('o053404, 16'o000000);
`MEM('o053406, 16'o000000);
`MEM('o053410, 16'o000000);
`MEM('o053412, 16'o000000);
`MEM('o053414, 16'o000000);
`MEM('o053416, 16'o000000);
`MEM('o053420, 16'o000000);
`MEM('o053422, 16'o000000);
`MEM('o053424, 16'o000000);
`MEM('o053426, 16'o000000);
`MEM('o053430, 16'o000000);
`MEM('o053432, 16'o000000);
`MEM('o053434, 16'o000000);
`MEM('o053436, 16'o000000);
`MEM('o053440, 16'o000000);
`MEM('o053442, 16'o000000);
`MEM('o053444, 16'o000000);
`MEM('o053446, 16'o000000);
`MEM('o053450, 16'o000000);
`MEM('o053452, 16'o000000);
`MEM('o053454, 16'o000000);
`MEM('o053456, 16'o000000);
`MEM('o053460, 16'o000000);
`MEM('o053462, 16'o000000);
`MEM('o053464, 16'o000000);
`MEM('o053466, 16'o000000);
`MEM('o053470, 16'o000000);
`MEM('o053472, 16'o000000);
`MEM('o053474, 16'o000000);
`MEM('o053476, 16'o000000);
`MEM('o053500, 16'o000000);
`MEM('o053502, 16'o000000);
`MEM('o053504, 16'o000000);
`MEM('o053506, 16'o000000);
`MEM('o053510, 16'o000000);
`MEM('o053512, 16'o000000);
`MEM('o053514, 16'o000000);
`MEM('o053516, 16'o000000);
`MEM('o053520, 16'o000000);
`MEM('o053522, 16'o000000);
`MEM('o053524, 16'o000000);
`MEM('o053526, 16'o000000);
`MEM('o053530, 16'o000000);
`MEM('o053532, 16'o000000);
`MEM('o053534, 16'o000000);
`MEM('o053536, 16'o000000);
`MEM('o053540, 16'o000000);
`MEM('o053542, 16'o000000);
`MEM('o053544, 16'o000000);
`MEM('o053546, 16'o000000);
`MEM('o053550, 16'o000000);
`MEM('o053552, 16'o000000);
`MEM('o053554, 16'o000000);
`MEM('o053556, 16'o000000);
`MEM('o053560, 16'o000000);
`MEM('o053562, 16'o000000);
`MEM('o053564, 16'o000000);
`MEM('o053566, 16'o000000);
`MEM('o053570, 16'o000000);
`MEM('o053572, 16'o000000);
`MEM('o053574, 16'o000000);
`MEM('o053576, 16'o000000);
`MEM('o053600, 16'o000000);
`MEM('o053602, 16'o000000);
`MEM('o053604, 16'o000000);
`MEM('o053606, 16'o000000);
`MEM('o053610, 16'o000000);
`MEM('o053612, 16'o000000);
`MEM('o053614, 16'o000000);
`MEM('o053616, 16'o000000);
`MEM('o053620, 16'o000000);
`MEM('o053622, 16'o000000);
`MEM('o053624, 16'o000000);
`MEM('o053626, 16'o000000);
`MEM('o053630, 16'o000000);
`MEM('o053632, 16'o000000);
`MEM('o053634, 16'o000000);
`MEM('o053636, 16'o000000);
`MEM('o053640, 16'o000000);
`MEM('o053642, 16'o000000);
`MEM('o053644, 16'o000000);
`MEM('o053646, 16'o000000);
`MEM('o053650, 16'o000000);
`MEM('o053652, 16'o000000);
`MEM('o053654, 16'o000000);
`MEM('o053656, 16'o000000);
`MEM('o053660, 16'o000000);
`MEM('o053662, 16'o000000);
`MEM('o053664, 16'o000000);
`MEM('o053666, 16'o000000);
`MEM('o053670, 16'o000000);
`MEM('o053672, 16'o000000);
`MEM('o053674, 16'o000000);
`MEM('o053676, 16'o000000);
`MEM('o053700, 16'o000000);
`MEM('o053702, 16'o000000);
`MEM('o053704, 16'o000000);
`MEM('o053706, 16'o000000);
`MEM('o053710, 16'o000000);
`MEM('o053712, 16'o000000);
`MEM('o053714, 16'o000000);
`MEM('o053716, 16'o000000);
`MEM('o053720, 16'o000000);
`MEM('o053722, 16'o000000);
`MEM('o053724, 16'o000000);
`MEM('o053726, 16'o000000);
`MEM('o053730, 16'o000000);
`MEM('o053732, 16'o000000);
`MEM('o053734, 16'o000000);
`MEM('o053736, 16'o000000);
`MEM('o053740, 16'o000000);
`MEM('o053742, 16'o000000);
`MEM('o053744, 16'o000000);
`MEM('o053746, 16'o000000);
`MEM('o053750, 16'o000000);
`MEM('o053752, 16'o000000);
`MEM('o053754, 16'o000000);
`MEM('o053756, 16'o000000);
`MEM('o053760, 16'o000000);
`MEM('o053762, 16'o000000);
`MEM('o053764, 16'o000000);
`MEM('o053766, 16'o000000);
`MEM('o053770, 16'o000000);
`MEM('o053772, 16'o000000);
`MEM('o053774, 16'o000000);
`MEM('o053776, 16'o000000);
`MEM('o054000, 16'o000000);
`MEM('o054002, 16'o000000);
`MEM('o054004, 16'o000000);
`MEM('o054006, 16'o000000);
`MEM('o054010, 16'o000000);
`MEM('o054012, 16'o000000);
`MEM('o054014, 16'o000000);
`MEM('o054016, 16'o000000);
`MEM('o054020, 16'o000000);
`MEM('o054022, 16'o000000);
`MEM('o054024, 16'o000000);
`MEM('o054026, 16'o000000);
`MEM('o054030, 16'o000000);
`MEM('o054032, 16'o000000);
`MEM('o054034, 16'o000000);
`MEM('o054036, 16'o000000);
`MEM('o054040, 16'o000000);
`MEM('o054042, 16'o000000);
`MEM('o054044, 16'o000000);
`MEM('o054046, 16'o000000);
`MEM('o054050, 16'o000000);
`MEM('o054052, 16'o000000);
`MEM('o054054, 16'o000000);
`MEM('o054056, 16'o000000);
`MEM('o054060, 16'o000000);
`MEM('o054062, 16'o000000);
`MEM('o054064, 16'o000000);
`MEM('o054066, 16'o000000);
`MEM('o054070, 16'o000000);
`MEM('o054072, 16'o000000);
`MEM('o054074, 16'o000000);
`MEM('o054076, 16'o000000);
`MEM('o054100, 16'o000000);
`MEM('o054102, 16'o000000);
`MEM('o054104, 16'o000000);
`MEM('o054106, 16'o000000);
`MEM('o054110, 16'o000000);
`MEM('o054112, 16'o000000);
`MEM('o054114, 16'o000000);
`MEM('o054116, 16'o000000);
`MEM('o054120, 16'o000000);
`MEM('o054122, 16'o000000);
`MEM('o054124, 16'o000000);
`MEM('o054126, 16'o000000);
`MEM('o054130, 16'o000000);
`MEM('o054132, 16'o000000);
`MEM('o054134, 16'o000000);
`MEM('o054136, 16'o000000);
`MEM('o054140, 16'o000000);
`MEM('o054142, 16'o000000);
`MEM('o054144, 16'o000000);
`MEM('o054146, 16'o000000);
`MEM('o054150, 16'o000000);
`MEM('o054152, 16'o000000);
`MEM('o054154, 16'o000000);
`MEM('o054156, 16'o000000);
`MEM('o054160, 16'o000000);
`MEM('o054162, 16'o000000);
`MEM('o054164, 16'o000000);
`MEM('o054166, 16'o000000);
`MEM('o054170, 16'o000000);
`MEM('o054172, 16'o000000);
`MEM('o054174, 16'o000000);
`MEM('o054176, 16'o000000);
`MEM('o054200, 16'o000000);
`MEM('o054202, 16'o000000);
`MEM('o054204, 16'o000000);
`MEM('o054206, 16'o000000);
`MEM('o054210, 16'o000000);
`MEM('o054212, 16'o000000);
`MEM('o054214, 16'o000000);
`MEM('o054216, 16'o000000);
`MEM('o054220, 16'o000000);
`MEM('o054222, 16'o000000);
`MEM('o054224, 16'o000000);
`MEM('o054226, 16'o000000);
`MEM('o054230, 16'o000000);
`MEM('o054232, 16'o000000);
`MEM('o054234, 16'o000000);
`MEM('o054236, 16'o000000);
`MEM('o054240, 16'o000000);
`MEM('o054242, 16'o000000);
`MEM('o054244, 16'o000000);
`MEM('o054246, 16'o000000);
`MEM('o054250, 16'o000000);
`MEM('o054252, 16'o000000);
`MEM('o054254, 16'o000000);
`MEM('o054256, 16'o000000);
`MEM('o054260, 16'o000000);
`MEM('o054262, 16'o000000);
`MEM('o054264, 16'o000000);
`MEM('o054266, 16'o000000);
`MEM('o054270, 16'o000000);
`MEM('o054272, 16'o000000);
`MEM('o054274, 16'o000000);
`MEM('o054276, 16'o000000);
`MEM('o054300, 16'o000000);
`MEM('o054302, 16'o000000);
`MEM('o054304, 16'o000000);
`MEM('o054306, 16'o000000);
`MEM('o054310, 16'o000000);
`MEM('o054312, 16'o000000);
`MEM('o054314, 16'o000000);
`MEM('o054316, 16'o000000);
`MEM('o054320, 16'o000000);
`MEM('o054322, 16'o000000);
`MEM('o054324, 16'o000000);
`MEM('o054326, 16'o000000);
`MEM('o054330, 16'o000000);
`MEM('o054332, 16'o000000);
`MEM('o054334, 16'o000000);
`MEM('o054336, 16'o000000);
`MEM('o054340, 16'o000000);
`MEM('o054342, 16'o000000);
`MEM('o054344, 16'o000000);
`MEM('o054346, 16'o000000);
`MEM('o054350, 16'o000000);
`MEM('o054352, 16'o000000);
`MEM('o054354, 16'o000000);
`MEM('o054356, 16'o000000);
`MEM('o054360, 16'o000000);
`MEM('o054362, 16'o000000);
`MEM('o054364, 16'o000000);
`MEM('o054366, 16'o000000);
`MEM('o054370, 16'o000000);
`MEM('o054372, 16'o000000);
`MEM('o054374, 16'o000000);
`MEM('o054376, 16'o000000);
`MEM('o054400, 16'o000000);
`MEM('o054402, 16'o000000);
`MEM('o054404, 16'o000000);
`MEM('o054406, 16'o000000);
`MEM('o054410, 16'o000000);
`MEM('o054412, 16'o000000);
`MEM('o054414, 16'o000000);
`MEM('o054416, 16'o000000);
`MEM('o054420, 16'o000000);
`MEM('o054422, 16'o000000);
`MEM('o054424, 16'o000000);
`MEM('o054426, 16'o000000);
`MEM('o054430, 16'o000000);
`MEM('o054432, 16'o000000);
`MEM('o054434, 16'o000000);
`MEM('o054436, 16'o000000);
`MEM('o054440, 16'o000000);
`MEM('o054442, 16'o000000);
`MEM('o054444, 16'o000000);
`MEM('o054446, 16'o000000);
`MEM('o054450, 16'o000000);
`MEM('o054452, 16'o000000);
`MEM('o054454, 16'o000000);
`MEM('o054456, 16'o000000);
`MEM('o054460, 16'o000000);
`MEM('o054462, 16'o000000);
`MEM('o054464, 16'o000000);
`MEM('o054466, 16'o000000);
`MEM('o054470, 16'o000000);
`MEM('o054472, 16'o000000);
`MEM('o054474, 16'o000000);
`MEM('o054476, 16'o000000);
`MEM('o054500, 16'o000000);
`MEM('o054502, 16'o000000);
`MEM('o054504, 16'o000000);
`MEM('o054506, 16'o000000);
`MEM('o054510, 16'o000000);
`MEM('o054512, 16'o000000);
`MEM('o054514, 16'o000000);
`MEM('o054516, 16'o000000);
`MEM('o054520, 16'o000000);
`MEM('o054522, 16'o000000);
`MEM('o054524, 16'o000000);
`MEM('o054526, 16'o000000);
`MEM('o054530, 16'o000000);
`MEM('o054532, 16'o000000);
`MEM('o054534, 16'o000000);
`MEM('o054536, 16'o000000);
`MEM('o054540, 16'o000000);
`MEM('o054542, 16'o000000);
`MEM('o054544, 16'o000000);
`MEM('o054546, 16'o000000);
`MEM('o054550, 16'o000000);
`MEM('o054552, 16'o000000);
`MEM('o054554, 16'o000000);
`MEM('o054556, 16'o000000);
`MEM('o054560, 16'o000000);
`MEM('o054562, 16'o000000);
`MEM('o054564, 16'o000000);
`MEM('o054566, 16'o000000);
`MEM('o054570, 16'o000000);
`MEM('o054572, 16'o000000);
`MEM('o054574, 16'o000000);
`MEM('o054576, 16'o000000);
`MEM('o054600, 16'o000000);
`MEM('o054602, 16'o000000);
`MEM('o054604, 16'o000000);
`MEM('o054606, 16'o000000);
`MEM('o054610, 16'o000000);
`MEM('o054612, 16'o000000);
`MEM('o054614, 16'o000000);
`MEM('o054616, 16'o000000);
`MEM('o054620, 16'o000000);
`MEM('o054622, 16'o000000);
`MEM('o054624, 16'o000000);
`MEM('o054626, 16'o000000);
`MEM('o054630, 16'o000000);
`MEM('o054632, 16'o000000);
`MEM('o054634, 16'o000000);
`MEM('o054636, 16'o000000);
`MEM('o054640, 16'o000000);
`MEM('o054642, 16'o000000);
`MEM('o054644, 16'o000000);
`MEM('o054646, 16'o000000);
`MEM('o054650, 16'o000000);
`MEM('o054652, 16'o000000);
`MEM('o054654, 16'o000000);
`MEM('o054656, 16'o000000);
`MEM('o054660, 16'o000000);
`MEM('o054662, 16'o000000);
`MEM('o054664, 16'o000000);
`MEM('o054666, 16'o000000);
`MEM('o054670, 16'o000000);
`MEM('o054672, 16'o000000);
`MEM('o054674, 16'o000000);
`MEM('o054676, 16'o000000);
`MEM('o054700, 16'o000000);
`MEM('o054702, 16'o000000);
`MEM('o054704, 16'o000000);
`MEM('o054706, 16'o000000);
`MEM('o054710, 16'o000000);
`MEM('o054712, 16'o000000);
`MEM('o054714, 16'o000000);
`MEM('o054716, 16'o000000);
`MEM('o054720, 16'o000000);
`MEM('o054722, 16'o000000);
`MEM('o054724, 16'o000000);
`MEM('o054726, 16'o000000);
`MEM('o054730, 16'o000000);
`MEM('o054732, 16'o000000);
`MEM('o054734, 16'o000000);
`MEM('o054736, 16'o000000);
`MEM('o054740, 16'o000000);
`MEM('o054742, 16'o000000);
`MEM('o054744, 16'o000000);
`MEM('o054746, 16'o000000);
`MEM('o054750, 16'o000000);
`MEM('o054752, 16'o000000);
`MEM('o054754, 16'o000000);
`MEM('o054756, 16'o000000);
`MEM('o054760, 16'o000000);
`MEM('o054762, 16'o000000);
`MEM('o054764, 16'o000000);
`MEM('o054766, 16'o000000);
`MEM('o054770, 16'o000000);
`MEM('o054772, 16'o000000);
`MEM('o054774, 16'o000000);
`MEM('o054776, 16'o000000);
`MEM('o055000, 16'o000000);
`MEM('o055002, 16'o000000);
`MEM('o055004, 16'o000000);
`MEM('o055006, 16'o000000);
`MEM('o055010, 16'o000000);
`MEM('o055012, 16'o000000);
`MEM('o055014, 16'o000000);
`MEM('o055016, 16'o000000);
`MEM('o055020, 16'o000000);
`MEM('o055022, 16'o000000);
`MEM('o055024, 16'o000000);
`MEM('o055026, 16'o000000);
`MEM('o055030, 16'o000000);
`MEM('o055032, 16'o000000);
`MEM('o055034, 16'o000000);
`MEM('o055036, 16'o000000);
`MEM('o055040, 16'o000000);
`MEM('o055042, 16'o000000);
`MEM('o055044, 16'o000000);
`MEM('o055046, 16'o000000);
`MEM('o055050, 16'o000000);
`MEM('o055052, 16'o000000);
`MEM('o055054, 16'o000000);
`MEM('o055056, 16'o000000);
`MEM('o055060, 16'o000000);
`MEM('o055062, 16'o000000);
`MEM('o055064, 16'o000000);
`MEM('o055066, 16'o000000);
`MEM('o055070, 16'o000000);
`MEM('o055072, 16'o000000);
`MEM('o055074, 16'o000000);
`MEM('o055076, 16'o000000);
`MEM('o055100, 16'o000000);
`MEM('o055102, 16'o000000);
`MEM('o055104, 16'o000000);
`MEM('o055106, 16'o000000);
`MEM('o055110, 16'o000000);
`MEM('o055112, 16'o000000);
`MEM('o055114, 16'o000000);
`MEM('o055116, 16'o000000);
`MEM('o055120, 16'o000000);
`MEM('o055122, 16'o000000);
`MEM('o055124, 16'o000000);
`MEM('o055126, 16'o000000);
`MEM('o055130, 16'o000000);
`MEM('o055132, 16'o000000);
`MEM('o055134, 16'o000000);
`MEM('o055136, 16'o000000);
`MEM('o055140, 16'o000000);
`MEM('o055142, 16'o000000);
`MEM('o055144, 16'o000000);
`MEM('o055146, 16'o000000);
`MEM('o055150, 16'o000000);
`MEM('o055152, 16'o000000);
`MEM('o055154, 16'o000000);
`MEM('o055156, 16'o000000);
`MEM('o055160, 16'o000000);
`MEM('o055162, 16'o000000);
`MEM('o055164, 16'o000000);
`MEM('o055166, 16'o000000);
`MEM('o055170, 16'o000000);
`MEM('o055172, 16'o000000);
`MEM('o055174, 16'o000000);
`MEM('o055176, 16'o000000);
`MEM('o055200, 16'o000000);
`MEM('o055202, 16'o000000);
`MEM('o055204, 16'o000000);
`MEM('o055206, 16'o000000);
`MEM('o055210, 16'o000000);
`MEM('o055212, 16'o000000);
`MEM('o055214, 16'o000000);
`MEM('o055216, 16'o000000);
`MEM('o055220, 16'o000000);
`MEM('o055222, 16'o000000);
`MEM('o055224, 16'o000000);
`MEM('o055226, 16'o000000);
`MEM('o055230, 16'o000000);
`MEM('o055232, 16'o000000);
`MEM('o055234, 16'o000000);
`MEM('o055236, 16'o000000);
`MEM('o055240, 16'o000000);
`MEM('o055242, 16'o000000);
`MEM('o055244, 16'o000000);
`MEM('o055246, 16'o000000);
`MEM('o055250, 16'o000000);
`MEM('o055252, 16'o000000);
`MEM('o055254, 16'o000000);
`MEM('o055256, 16'o000000);
`MEM('o055260, 16'o000000);
`MEM('o055262, 16'o000000);
`MEM('o055264, 16'o000000);
`MEM('o055266, 16'o000000);
`MEM('o055270, 16'o000000);
`MEM('o055272, 16'o000000);
`MEM('o055274, 16'o000000);
`MEM('o055276, 16'o000000);
`MEM('o055300, 16'o000000);
`MEM('o055302, 16'o000000);
`MEM('o055304, 16'o000000);
`MEM('o055306, 16'o000000);
`MEM('o055310, 16'o000000);
`MEM('o055312, 16'o000000);
`MEM('o055314, 16'o000000);
`MEM('o055316, 16'o000000);
`MEM('o055320, 16'o000000);
`MEM('o055322, 16'o000000);
`MEM('o055324, 16'o000000);
`MEM('o055326, 16'o000000);
`MEM('o055330, 16'o000000);
`MEM('o055332, 16'o000000);
`MEM('o055334, 16'o000000);
`MEM('o055336, 16'o000000);
`MEM('o055340, 16'o000000);
`MEM('o055342, 16'o000000);
`MEM('o055344, 16'o000000);
`MEM('o055346, 16'o000000);
`MEM('o055350, 16'o000000);
`MEM('o055352, 16'o000000);
`MEM('o055354, 16'o000000);
`MEM('o055356, 16'o000000);
`MEM('o055360, 16'o000000);
`MEM('o055362, 16'o000000);
`MEM('o055364, 16'o000000);
`MEM('o055366, 16'o000000);
`MEM('o055370, 16'o000000);
`MEM('o055372, 16'o000000);
`MEM('o055374, 16'o000000);
`MEM('o055376, 16'o000000);
`MEM('o055400, 16'o000000);
`MEM('o055402, 16'o000000);
`MEM('o055404, 16'o000000);
`MEM('o055406, 16'o000000);
`MEM('o055410, 16'o000000);
`MEM('o055412, 16'o000000);
`MEM('o055414, 16'o000000);
`MEM('o055416, 16'o000000);
`MEM('o055420, 16'o000000);
`MEM('o055422, 16'o000000);
`MEM('o055424, 16'o000000);
`MEM('o055426, 16'o000000);
`MEM('o055430, 16'o000000);
`MEM('o055432, 16'o000000);
`MEM('o055434, 16'o000000);
`MEM('o055436, 16'o000000);
`MEM('o055440, 16'o000000);
`MEM('o055442, 16'o000000);
`MEM('o055444, 16'o000000);
`MEM('o055446, 16'o000000);
`MEM('o055450, 16'o000000);
`MEM('o055452, 16'o000000);
`MEM('o055454, 16'o000000);
`MEM('o055456, 16'o000000);
`MEM('o055460, 16'o000000);
`MEM('o055462, 16'o000000);
`MEM('o055464, 16'o000000);
`MEM('o055466, 16'o000000);
`MEM('o055470, 16'o000000);
`MEM('o055472, 16'o000000);
`MEM('o055474, 16'o000000);
`MEM('o055476, 16'o000000);
`MEM('o055500, 16'o000000);
`MEM('o055502, 16'o000000);
`MEM('o055504, 16'o000000);
`MEM('o055506, 16'o000000);
`MEM('o055510, 16'o000000);
`MEM('o055512, 16'o000000);
`MEM('o055514, 16'o000000);
`MEM('o055516, 16'o000000);
`MEM('o055520, 16'o000000);
`MEM('o055522, 16'o000000);
`MEM('o055524, 16'o000000);
`MEM('o055526, 16'o000000);
`MEM('o055530, 16'o000000);
`MEM('o055532, 16'o000000);
`MEM('o055534, 16'o000000);
`MEM('o055536, 16'o000000);
`MEM('o055540, 16'o000000);
`MEM('o055542, 16'o000000);
`MEM('o055544, 16'o000000);
`MEM('o055546, 16'o000000);
`MEM('o055550, 16'o000000);
`MEM('o055552, 16'o000000);
`MEM('o055554, 16'o000000);
`MEM('o055556, 16'o000000);
`MEM('o055560, 16'o000000);
`MEM('o055562, 16'o000000);
`MEM('o055564, 16'o000000);
`MEM('o055566, 16'o000000);
`MEM('o055570, 16'o000000);
`MEM('o055572, 16'o000000);
`MEM('o055574, 16'o000000);
`MEM('o055576, 16'o000000);
`MEM('o055600, 16'o000000);
`MEM('o055602, 16'o000000);
`MEM('o055604, 16'o000000);
`MEM('o055606, 16'o000000);
`MEM('o055610, 16'o000000);
`MEM('o055612, 16'o000000);
`MEM('o055614, 16'o000000);
`MEM('o055616, 16'o000000);
`MEM('o055620, 16'o000000);
`MEM('o055622, 16'o000000);
`MEM('o055624, 16'o000000);
`MEM('o055626, 16'o000000);
`MEM('o055630, 16'o000000);
`MEM('o055632, 16'o000000);
`MEM('o055634, 16'o000000);
`MEM('o055636, 16'o000000);
`MEM('o055640, 16'o000000);
`MEM('o055642, 16'o000000);
`MEM('o055644, 16'o000000);
`MEM('o055646, 16'o000000);
`MEM('o055650, 16'o000000);
`MEM('o055652, 16'o000000);
`MEM('o055654, 16'o000000);
`MEM('o055656, 16'o000000);
`MEM('o055660, 16'o000000);
`MEM('o055662, 16'o000000);
`MEM('o055664, 16'o000000);
`MEM('o055666, 16'o000000);
`MEM('o055670, 16'o000000);
`MEM('o055672, 16'o000000);
`MEM('o055674, 16'o000000);
`MEM('o055676, 16'o000000);
`MEM('o055700, 16'o000000);
`MEM('o055702, 16'o000000);
`MEM('o055704, 16'o000000);
`MEM('o055706, 16'o000000);
`MEM('o055710, 16'o000000);
`MEM('o055712, 16'o000000);
`MEM('o055714, 16'o000000);
`MEM('o055716, 16'o000000);
`MEM('o055720, 16'o000000);
`MEM('o055722, 16'o000000);
`MEM('o055724, 16'o000000);
`MEM('o055726, 16'o000000);
`MEM('o055730, 16'o000000);
`MEM('o055732, 16'o000000);
`MEM('o055734, 16'o000000);
`MEM('o055736, 16'o000000);
`MEM('o055740, 16'o000000);
`MEM('o055742, 16'o000000);
`MEM('o055744, 16'o000000);
`MEM('o055746, 16'o000000);
`MEM('o055750, 16'o000000);
`MEM('o055752, 16'o000000);
`MEM('o055754, 16'o000000);
`MEM('o055756, 16'o000000);
`MEM('o055760, 16'o000000);
`MEM('o055762, 16'o000000);
`MEM('o055764, 16'o000000);
`MEM('o055766, 16'o000000);
`MEM('o055770, 16'o000000);
`MEM('o055772, 16'o000000);
`MEM('o055774, 16'o000000);
`MEM('o055776, 16'o000000);
`MEM('o056000, 16'o000000);
`MEM('o056002, 16'o000000);
`MEM('o056004, 16'o000000);
`MEM('o056006, 16'o000000);
`MEM('o056010, 16'o000000);
`MEM('o056012, 16'o000000);
`MEM('o056014, 16'o000000);
`MEM('o056016, 16'o000000);
`MEM('o056020, 16'o000000);
`MEM('o056022, 16'o000000);
`MEM('o056024, 16'o000000);
`MEM('o056026, 16'o000000);
`MEM('o056030, 16'o000000);
`MEM('o056032, 16'o000000);
`MEM('o056034, 16'o000000);
`MEM('o056036, 16'o000000);
`MEM('o056040, 16'o000000);
`MEM('o056042, 16'o000000);
`MEM('o056044, 16'o000000);
`MEM('o056046, 16'o000000);
`MEM('o056050, 16'o000000);
`MEM('o056052, 16'o000000);
`MEM('o056054, 16'o000000);
`MEM('o056056, 16'o000000);
`MEM('o056060, 16'o000000);
`MEM('o056062, 16'o000000);
`MEM('o056064, 16'o000000);
`MEM('o056066, 16'o000000);
`MEM('o056070, 16'o000000);
`MEM('o056072, 16'o000000);
`MEM('o056074, 16'o000000);
`MEM('o056076, 16'o000000);
`MEM('o056100, 16'o000000);
`MEM('o056102, 16'o000000);
`MEM('o056104, 16'o000000);
`MEM('o056106, 16'o000000);
`MEM('o056110, 16'o000000);
`MEM('o056112, 16'o000000);
`MEM('o056114, 16'o000000);
`MEM('o056116, 16'o000000);
`MEM('o056120, 16'o000000);
`MEM('o056122, 16'o000000);
`MEM('o056124, 16'o000000);
`MEM('o056126, 16'o000000);
`MEM('o056130, 16'o000000);
`MEM('o056132, 16'o000000);
`MEM('o056134, 16'o000000);
`MEM('o056136, 16'o000000);
`MEM('o056140, 16'o000000);
`MEM('o056142, 16'o000000);
`MEM('o056144, 16'o000000);
`MEM('o056146, 16'o000000);
`MEM('o056150, 16'o000000);
`MEM('o056152, 16'o000000);
`MEM('o056154, 16'o000000);
`MEM('o056156, 16'o000000);
`MEM('o056160, 16'o000000);
`MEM('o056162, 16'o000000);
`MEM('o056164, 16'o000000);
`MEM('o056166, 16'o000000);
`MEM('o056170, 16'o000000);
`MEM('o056172, 16'o000000);
`MEM('o056174, 16'o000000);
`MEM('o056176, 16'o000000);
`MEM('o056200, 16'o000000);
`MEM('o056202, 16'o000000);
`MEM('o056204, 16'o000000);
`MEM('o056206, 16'o000000);
`MEM('o056210, 16'o000000);
`MEM('o056212, 16'o000000);
`MEM('o056214, 16'o000000);
`MEM('o056216, 16'o000000);
`MEM('o056220, 16'o000000);
`MEM('o056222, 16'o000000);
`MEM('o056224, 16'o000000);
`MEM('o056226, 16'o000000);
`MEM('o056230, 16'o000000);
`MEM('o056232, 16'o000000);
`MEM('o056234, 16'o000000);
`MEM('o056236, 16'o000000);
`MEM('o056240, 16'o000000);
`MEM('o056242, 16'o000000);
`MEM('o056244, 16'o000000);
`MEM('o056246, 16'o000000);
`MEM('o056250, 16'o000000);
`MEM('o056252, 16'o000000);
`MEM('o056254, 16'o000000);
`MEM('o056256, 16'o000000);
`MEM('o056260, 16'o000000);
`MEM('o056262, 16'o000000);
`MEM('o056264, 16'o000000);
`MEM('o056266, 16'o000000);
`MEM('o056270, 16'o000000);
`MEM('o056272, 16'o000000);
`MEM('o056274, 16'o000000);
`MEM('o056276, 16'o000000);
`MEM('o056300, 16'o000000);
`MEM('o056302, 16'o000000);
`MEM('o056304, 16'o000000);
`MEM('o056306, 16'o000000);
`MEM('o056310, 16'o000000);
`MEM('o056312, 16'o000000);
`MEM('o056314, 16'o000000);
`MEM('o056316, 16'o000000);
`MEM('o056320, 16'o000000);
`MEM('o056322, 16'o000000);
`MEM('o056324, 16'o000000);
`MEM('o056326, 16'o000000);
`MEM('o056330, 16'o000000);
`MEM('o056332, 16'o000000);
`MEM('o056334, 16'o000000);
`MEM('o056336, 16'o000000);
`MEM('o056340, 16'o000000);
`MEM('o056342, 16'o000000);
`MEM('o056344, 16'o000000);
`MEM('o056346, 16'o000000);
`MEM('o056350, 16'o000000);
`MEM('o056352, 16'o000000);
`MEM('o056354, 16'o000000);
`MEM('o056356, 16'o000000);
`MEM('o056360, 16'o000000);
`MEM('o056362, 16'o000000);
`MEM('o056364, 16'o000000);
`MEM('o056366, 16'o000000);
`MEM('o056370, 16'o000000);
`MEM('o056372, 16'o000000);
`MEM('o056374, 16'o000000);
`MEM('o056376, 16'o000000);
`MEM('o056400, 16'o000000);
`MEM('o056402, 16'o000000);
`MEM('o056404, 16'o000000);
`MEM('o056406, 16'o000000);
`MEM('o056410, 16'o000000);
`MEM('o056412, 16'o000000);
`MEM('o056414, 16'o000000);
`MEM('o056416, 16'o000000);
`MEM('o056420, 16'o000000);
`MEM('o056422, 16'o000000);
`MEM('o056424, 16'o000000);
`MEM('o056426, 16'o000000);
`MEM('o056430, 16'o000000);
`MEM('o056432, 16'o000000);
`MEM('o056434, 16'o000000);
`MEM('o056436, 16'o000000);
`MEM('o056440, 16'o000000);
`MEM('o056442, 16'o000000);
`MEM('o056444, 16'o000000);
`MEM('o056446, 16'o000000);
`MEM('o056450, 16'o000000);
`MEM('o056452, 16'o000000);
`MEM('o056454, 16'o000000);
`MEM('o056456, 16'o000000);
`MEM('o056460, 16'o000000);
`MEM('o056462, 16'o000000);
`MEM('o056464, 16'o000000);
`MEM('o056466, 16'o000000);
`MEM('o056470, 16'o000000);
`MEM('o056472, 16'o000000);
`MEM('o056474, 16'o000000);
`MEM('o056476, 16'o000000);
`MEM('o056500, 16'o000000);
`MEM('o056502, 16'o000000);
`MEM('o056504, 16'o000000);
`MEM('o056506, 16'o000000);
`MEM('o056510, 16'o000000);
`MEM('o056512, 16'o000000);
`MEM('o056514, 16'o000000);
`MEM('o056516, 16'o000000);
`MEM('o056520, 16'o000000);
`MEM('o056522, 16'o000000);
`MEM('o056524, 16'o000000);
`MEM('o056526, 16'o000000);
`MEM('o056530, 16'o000000);
`MEM('o056532, 16'o000000);
`MEM('o056534, 16'o000000);
`MEM('o056536, 16'o000000);
`MEM('o056540, 16'o000000);
`MEM('o056542, 16'o000000);
`MEM('o056544, 16'o000000);
`MEM('o056546, 16'o000000);
`MEM('o056550, 16'o000000);
`MEM('o056552, 16'o000000);
`MEM('o056554, 16'o000000);
`MEM('o056556, 16'o000000);
`MEM('o056560, 16'o000000);
`MEM('o056562, 16'o000000);
`MEM('o056564, 16'o000000);
`MEM('o056566, 16'o000000);
`MEM('o056570, 16'o000000);
`MEM('o056572, 16'o000000);
`MEM('o056574, 16'o000000);
`MEM('o056576, 16'o000000);
`MEM('o056600, 16'o000000);
`MEM('o056602, 16'o000000);
`MEM('o056604, 16'o000000);
`MEM('o056606, 16'o000000);
`MEM('o056610, 16'o000000);
`MEM('o056612, 16'o000000);
`MEM('o056614, 16'o000000);
`MEM('o056616, 16'o000000);
`MEM('o056620, 16'o000000);
`MEM('o056622, 16'o000000);
`MEM('o056624, 16'o000000);
`MEM('o056626, 16'o000000);
`MEM('o056630, 16'o000000);
`MEM('o056632, 16'o000000);
`MEM('o056634, 16'o000000);
`MEM('o056636, 16'o000000);
`MEM('o056640, 16'o000000);
`MEM('o056642, 16'o000000);
`MEM('o056644, 16'o000000);
`MEM('o056646, 16'o000000);
`MEM('o056650, 16'o000000);
`MEM('o056652, 16'o000000);
`MEM('o056654, 16'o000000);
`MEM('o056656, 16'o000000);
`MEM('o056660, 16'o000000);
`MEM('o056662, 16'o000000);
`MEM('o056664, 16'o000000);
`MEM('o056666, 16'o000000);
`MEM('o056670, 16'o000000);
`MEM('o056672, 16'o000000);
`MEM('o056674, 16'o000000);
`MEM('o056676, 16'o000000);
`MEM('o056700, 16'o000000);
`MEM('o056702, 16'o000000);
`MEM('o056704, 16'o000000);
`MEM('o056706, 16'o000000);
`MEM('o056710, 16'o000000);
`MEM('o056712, 16'o000000);
`MEM('o056714, 16'o000000);
`MEM('o056716, 16'o000000);
`MEM('o056720, 16'o000000);
`MEM('o056722, 16'o000000);
`MEM('o056724, 16'o000000);
`MEM('o056726, 16'o000000);
`MEM('o056730, 16'o000000);
`MEM('o056732, 16'o000000);
`MEM('o056734, 16'o000000);
`MEM('o056736, 16'o000000);
`MEM('o056740, 16'o000000);
`MEM('o056742, 16'o000000);
`MEM('o056744, 16'o000000);
`MEM('o056746, 16'o000000);
`MEM('o056750, 16'o000000);
`MEM('o056752, 16'o000000);
`MEM('o056754, 16'o000000);
`MEM('o056756, 16'o000000);
`MEM('o056760, 16'o000000);
`MEM('o056762, 16'o000000);
`MEM('o056764, 16'o000000);
`MEM('o056766, 16'o000000);
`MEM('o056770, 16'o000000);
`MEM('o056772, 16'o000000);
`MEM('o056774, 16'o000000);
`MEM('o056776, 16'o000000);
`MEM('o057000, 16'o000000);
`MEM('o057002, 16'o000000);
`MEM('o057004, 16'o000000);
`MEM('o057006, 16'o000000);
`MEM('o057010, 16'o000000);
`MEM('o057012, 16'o000000);
`MEM('o057014, 16'o000000);
`MEM('o057016, 16'o000000);
`MEM('o057020, 16'o000000);
`MEM('o057022, 16'o000000);
`MEM('o057024, 16'o000000);
`MEM('o057026, 16'o000000);
`MEM('o057030, 16'o000000);
`MEM('o057032, 16'o000000);
`MEM('o057034, 16'o000000);
`MEM('o057036, 16'o000000);
`MEM('o057040, 16'o000000);
`MEM('o057042, 16'o000000);
`MEM('o057044, 16'o000000);
`MEM('o057046, 16'o000000);
`MEM('o057050, 16'o000000);
`MEM('o057052, 16'o000000);
`MEM('o057054, 16'o000000);
`MEM('o057056, 16'o000000);
`MEM('o057060, 16'o000000);
`MEM('o057062, 16'o000000);
`MEM('o057064, 16'o000000);
`MEM('o057066, 16'o000000);
`MEM('o057070, 16'o000000);
`MEM('o057072, 16'o000000);
`MEM('o057074, 16'o000000);
`MEM('o057076, 16'o000000);
`MEM('o057100, 16'o000000);
`MEM('o057102, 16'o000000);
`MEM('o057104, 16'o000000);
`MEM('o057106, 16'o000000);
`MEM('o057110, 16'o000000);
`MEM('o057112, 16'o000000);
`MEM('o057114, 16'o000000);
`MEM('o057116, 16'o000000);
`MEM('o057120, 16'o000000);
`MEM('o057122, 16'o000000);
`MEM('o057124, 16'o000000);
`MEM('o057126, 16'o000000);
`MEM('o057130, 16'o000000);
`MEM('o057132, 16'o000000);
`MEM('o057134, 16'o000000);
`MEM('o057136, 16'o000000);
`MEM('o057140, 16'o000000);
`MEM('o057142, 16'o000000);
`MEM('o057144, 16'o000000);
`MEM('o057146, 16'o000000);
`MEM('o057150, 16'o000000);
`MEM('o057152, 16'o000000);
`MEM('o057154, 16'o000000);
`MEM('o057156, 16'o000000);
`MEM('o057160, 16'o000000);
`MEM('o057162, 16'o000000);
`MEM('o057164, 16'o000000);
`MEM('o057166, 16'o000000);
`MEM('o057170, 16'o000000);
`MEM('o057172, 16'o000000);
`MEM('o057174, 16'o000000);
`MEM('o057176, 16'o000000);
`MEM('o057200, 16'o000000);
`MEM('o057202, 16'o000000);
`MEM('o057204, 16'o000000);
`MEM('o057206, 16'o000000);
`MEM('o057210, 16'o000000);
`MEM('o057212, 16'o000000);
`MEM('o057214, 16'o000000);
`MEM('o057216, 16'o000000);
`MEM('o057220, 16'o000000);
`MEM('o057222, 16'o000000);
`MEM('o057224, 16'o000000);
`MEM('o057226, 16'o000000);
`MEM('o057230, 16'o000000);
`MEM('o057232, 16'o000000);
`MEM('o057234, 16'o000000);
`MEM('o057236, 16'o000000);
`MEM('o057240, 16'o000000);
`MEM('o057242, 16'o000000);
`MEM('o057244, 16'o000000);
`MEM('o057246, 16'o000000);
`MEM('o057250, 16'o000000);
`MEM('o057252, 16'o000000);
`MEM('o057254, 16'o000000);
`MEM('o057256, 16'o000000);
`MEM('o057260, 16'o000000);
`MEM('o057262, 16'o000000);
`MEM('o057264, 16'o000000);
`MEM('o057266, 16'o000000);
`MEM('o057270, 16'o000000);
`MEM('o057272, 16'o000000);
`MEM('o057274, 16'o000000);
`MEM('o057276, 16'o000000);
`MEM('o057300, 16'o000000);
`MEM('o057302, 16'o000000);
`MEM('o057304, 16'o000000);
`MEM('o057306, 16'o000000);
`MEM('o057310, 16'o000000);
`MEM('o057312, 16'o000000);
`MEM('o057314, 16'o000000);
`MEM('o057316, 16'o000000);
`MEM('o057320, 16'o000000);
`MEM('o057322, 16'o000000);
`MEM('o057324, 16'o000000);
`MEM('o057326, 16'o000000);
`MEM('o057330, 16'o000000);
`MEM('o057332, 16'o000000);
`MEM('o057334, 16'o000000);
`MEM('o057336, 16'o000000);
`MEM('o057340, 16'o000000);
`MEM('o057342, 16'o000000);
`MEM('o057344, 16'o000000);
`MEM('o057346, 16'o000000);
`MEM('o057350, 16'o000000);
`MEM('o057352, 16'o000000);
`MEM('o057354, 16'o000000);
`MEM('o057356, 16'o000000);
`MEM('o057360, 16'o000000);
`MEM('o057362, 16'o000000);
`MEM('o057364, 16'o000000);
`MEM('o057366, 16'o000000);
`MEM('o057370, 16'o000000);
`MEM('o057372, 16'o000000);
`MEM('o057374, 16'o000000);
`MEM('o057376, 16'o000000);
`MEM('o057400, 16'o000000);
`MEM('o057402, 16'o000000);
`MEM('o057404, 16'o000000);
`MEM('o057406, 16'o000000);
`MEM('o057410, 16'o000000);
`MEM('o057412, 16'o000000);
`MEM('o057414, 16'o000000);
`MEM('o057416, 16'o000000);
`MEM('o057420, 16'o000000);
`MEM('o057422, 16'o000000);
`MEM('o057424, 16'o000000);
`MEM('o057426, 16'o000000);
`MEM('o057430, 16'o000000);
`MEM('o057432, 16'o000000);
`MEM('o057434, 16'o000000);
`MEM('o057436, 16'o000000);
`MEM('o057440, 16'o000000);
`MEM('o057442, 16'o000000);
`MEM('o057444, 16'o000000);
`MEM('o057446, 16'o000000);
`MEM('o057450, 16'o000000);
`MEM('o057452, 16'o000000);
`MEM('o057454, 16'o000000);
`MEM('o057456, 16'o000000);
`MEM('o057460, 16'o000000);
`MEM('o057462, 16'o000000);
`MEM('o057464, 16'o000000);
`MEM('o057466, 16'o000000);
`MEM('o057470, 16'o000000);
`MEM('o057472, 16'o000000);
`MEM('o057474, 16'o000000);
`MEM('o057476, 16'o000000);
`MEM('o057500, 16'o000000);
`MEM('o057502, 16'o000000);
`MEM('o057504, 16'o000000);
`MEM('o057506, 16'o000000);
`MEM('o057510, 16'o000000);
`MEM('o057512, 16'o000000);
`MEM('o057514, 16'o000000);
`MEM('o057516, 16'o000000);
`MEM('o057520, 16'o000000);
`MEM('o057522, 16'o000000);
`MEM('o057524, 16'o000000);
`MEM('o057526, 16'o000000);
`MEM('o057530, 16'o000000);
`MEM('o057532, 16'o000000);
`MEM('o057534, 16'o000000);
`MEM('o057536, 16'o000000);
`MEM('o057540, 16'o000000);
`MEM('o057542, 16'o000000);
`MEM('o057544, 16'o000000);
`MEM('o057546, 16'o000000);
`MEM('o057550, 16'o000000);
`MEM('o057552, 16'o000000);
`MEM('o057554, 16'o000000);
`MEM('o057556, 16'o000000);
`MEM('o057560, 16'o000000);
`MEM('o057562, 16'o000000);
`MEM('o057564, 16'o000000);
`MEM('o057566, 16'o000000);
`MEM('o057570, 16'o000000);
`MEM('o057572, 16'o000000);
`MEM('o057574, 16'o000000);
`MEM('o057576, 16'o000000);
`MEM('o057600, 16'o000000);
`MEM('o057602, 16'o000000);
`MEM('o057604, 16'o000000);
`MEM('o057606, 16'o000000);
`MEM('o057610, 16'o000000);
`MEM('o057612, 16'o000000);
`MEM('o057614, 16'o000000);
`MEM('o057616, 16'o000000);
`MEM('o057620, 16'o000000);
`MEM('o057622, 16'o000000);
`MEM('o057624, 16'o000000);
`MEM('o057626, 16'o000000);
`MEM('o057630, 16'o000000);
`MEM('o057632, 16'o000000);
`MEM('o057634, 16'o000000);
`MEM('o057636, 16'o000000);
`MEM('o057640, 16'o000000);
`MEM('o057642, 16'o000000);
`MEM('o057644, 16'o000000);
`MEM('o057646, 16'o000000);
`MEM('o057650, 16'o000000);
`MEM('o057652, 16'o000000);
`MEM('o057654, 16'o000000);
`MEM('o057656, 16'o000000);
`MEM('o057660, 16'o000000);
`MEM('o057662, 16'o000000);
`MEM('o057664, 16'o000000);
`MEM('o057666, 16'o000000);
`MEM('o057670, 16'o000000);
`MEM('o057672, 16'o000000);
`MEM('o057674, 16'o000000);
`MEM('o057676, 16'o000000);
`MEM('o057700, 16'o000000);
`MEM('o057702, 16'o000000);
`MEM('o057704, 16'o000000);
`MEM('o057706, 16'o000000);
`MEM('o057710, 16'o000000);
`MEM('o057712, 16'o000000);
`MEM('o057714, 16'o000000);
`MEM('o057716, 16'o000000);
`MEM('o057720, 16'o000000);
`MEM('o057722, 16'o000000);
`MEM('o057724, 16'o000000);
`MEM('o057726, 16'o000000);
`MEM('o057730, 16'o000000);
`MEM('o057732, 16'o000000);
`MEM('o057734, 16'o000000);
`MEM('o057736, 16'o000000);
`MEM('o057740, 16'o000000);
`MEM('o057742, 16'o000000);
`MEM('o057744, 16'o000000);
`MEM('o057746, 16'o000000);
`MEM('o057750, 16'o000000);
`MEM('o057752, 16'o000000);
`MEM('o057754, 16'o000000);
`MEM('o057756, 16'o000000);
`MEM('o057760, 16'o000000);
`MEM('o057762, 16'o000000);
`MEM('o057764, 16'o000000);
`MEM('o057766, 16'o000000);
`MEM('o057770, 16'o000000);
`MEM('o057772, 16'o000000);
`MEM('o057774, 16'o000000);
`MEM('o057776, 16'o000000);
`MEM('o060000, 16'o000000);
`MEM('o060002, 16'o000000);
`MEM('o060004, 16'o000000);
`MEM('o060006, 16'o000000);
`MEM('o060010, 16'o000000);
`MEM('o060012, 16'o000000);
`MEM('o060014, 16'o000000);
`MEM('o060016, 16'o000000);
`MEM('o060020, 16'o000000);
`MEM('o060022, 16'o000000);
`MEM('o060024, 16'o000000);
`MEM('o060026, 16'o000000);
`MEM('o060030, 16'o000000);
`MEM('o060032, 16'o000000);
`MEM('o060034, 16'o000000);
`MEM('o060036, 16'o000000);
`MEM('o060040, 16'o000000);
`MEM('o060042, 16'o000000);
`MEM('o060044, 16'o000000);
`MEM('o060046, 16'o000000);
`MEM('o060050, 16'o000000);
`MEM('o060052, 16'o000000);
`MEM('o060054, 16'o000000);
`MEM('o060056, 16'o000000);
`MEM('o060060, 16'o000000);
`MEM('o060062, 16'o000000);
`MEM('o060064, 16'o000000);
`MEM('o060066, 16'o000000);
`MEM('o060070, 16'o000000);
`MEM('o060072, 16'o000000);
`MEM('o060074, 16'o000000);
`MEM('o060076, 16'o000000);
`MEM('o060100, 16'o000000);
`MEM('o060102, 16'o000000);
`MEM('o060104, 16'o000000);
`MEM('o060106, 16'o000000);
`MEM('o060110, 16'o000000);
`MEM('o060112, 16'o000000);
`MEM('o060114, 16'o000000);
`MEM('o060116, 16'o000000);
`MEM('o060120, 16'o000000);
`MEM('o060122, 16'o000000);
`MEM('o060124, 16'o000000);
`MEM('o060126, 16'o000000);
`MEM('o060130, 16'o000000);
`MEM('o060132, 16'o000000);
`MEM('o060134, 16'o000000);
`MEM('o060136, 16'o000000);
`MEM('o060140, 16'o000000);
`MEM('o060142, 16'o000000);
`MEM('o060144, 16'o000000);
`MEM('o060146, 16'o000000);
`MEM('o060150, 16'o000000);
`MEM('o060152, 16'o000000);
`MEM('o060154, 16'o000000);
`MEM('o060156, 16'o000000);
`MEM('o060160, 16'o000000);
`MEM('o060162, 16'o000000);
`MEM('o060164, 16'o000000);
`MEM('o060166, 16'o000000);
`MEM('o060170, 16'o000000);
`MEM('o060172, 16'o000000);
`MEM('o060174, 16'o000000);
`MEM('o060176, 16'o000000);
`MEM('o060200, 16'o000000);
`MEM('o060202, 16'o000000);
`MEM('o060204, 16'o000000);
`MEM('o060206, 16'o000000);
`MEM('o060210, 16'o000000);
`MEM('o060212, 16'o000000);
`MEM('o060214, 16'o000000);
`MEM('o060216, 16'o000000);
`MEM('o060220, 16'o000000);
`MEM('o060222, 16'o000000);
`MEM('o060224, 16'o000000);
`MEM('o060226, 16'o000000);
`MEM('o060230, 16'o000000);
`MEM('o060232, 16'o000000);
`MEM('o060234, 16'o000000);
`MEM('o060236, 16'o000000);
`MEM('o060240, 16'o000000);
`MEM('o060242, 16'o000000);
`MEM('o060244, 16'o000000);
`MEM('o060246, 16'o000000);
`MEM('o060250, 16'o000000);
`MEM('o060252, 16'o000000);
`MEM('o060254, 16'o000000);
`MEM('o060256, 16'o000000);
`MEM('o060260, 16'o000000);
`MEM('o060262, 16'o000000);
`MEM('o060264, 16'o000000);
`MEM('o060266, 16'o000000);
`MEM('o060270, 16'o000000);
`MEM('o060272, 16'o000000);
`MEM('o060274, 16'o000000);
`MEM('o060276, 16'o000000);
`MEM('o060300, 16'o000000);
`MEM('o060302, 16'o000000);
`MEM('o060304, 16'o000000);
`MEM('o060306, 16'o000000);
`MEM('o060310, 16'o000000);
`MEM('o060312, 16'o000000);
`MEM('o060314, 16'o000000);
`MEM('o060316, 16'o000000);
`MEM('o060320, 16'o000000);
`MEM('o060322, 16'o000000);
`MEM('o060324, 16'o000000);
`MEM('o060326, 16'o000000);
`MEM('o060330, 16'o000000);
`MEM('o060332, 16'o000000);
`MEM('o060334, 16'o000000);
`MEM('o060336, 16'o000000);
`MEM('o060340, 16'o000000);
`MEM('o060342, 16'o000000);
`MEM('o060344, 16'o000000);
`MEM('o060346, 16'o000000);
`MEM('o060350, 16'o000000);
`MEM('o060352, 16'o000000);
`MEM('o060354, 16'o000000);
`MEM('o060356, 16'o000000);
`MEM('o060360, 16'o000000);
`MEM('o060362, 16'o000000);
`MEM('o060364, 16'o000000);
`MEM('o060366, 16'o000000);
`MEM('o060370, 16'o000000);
`MEM('o060372, 16'o000000);
`MEM('o060374, 16'o000000);
`MEM('o060376, 16'o000000);
`MEM('o060400, 16'o000000);
`MEM('o060402, 16'o000000);
`MEM('o060404, 16'o000000);
`MEM('o060406, 16'o000000);
`MEM('o060410, 16'o000000);
`MEM('o060412, 16'o000000);
`MEM('o060414, 16'o000000);
`MEM('o060416, 16'o000000);
`MEM('o060420, 16'o000000);
`MEM('o060422, 16'o000000);
`MEM('o060424, 16'o000000);
`MEM('o060426, 16'o000000);
`MEM('o060430, 16'o000000);
`MEM('o060432, 16'o000000);
`MEM('o060434, 16'o000000);
`MEM('o060436, 16'o000000);
`MEM('o060440, 16'o000000);
`MEM('o060442, 16'o000000);
`MEM('o060444, 16'o000000);
`MEM('o060446, 16'o000000);
`MEM('o060450, 16'o000000);
`MEM('o060452, 16'o000000);
`MEM('o060454, 16'o000000);
`MEM('o060456, 16'o000000);
`MEM('o060460, 16'o000000);
`MEM('o060462, 16'o000000);
`MEM('o060464, 16'o000000);
`MEM('o060466, 16'o000000);
`MEM('o060470, 16'o000000);
`MEM('o060472, 16'o000000);
`MEM('o060474, 16'o000000);
`MEM('o060476, 16'o000000);
`MEM('o060500, 16'o000000);
`MEM('o060502, 16'o000000);
`MEM('o060504, 16'o000000);
`MEM('o060506, 16'o000000);
`MEM('o060510, 16'o000000);
`MEM('o060512, 16'o000000);
`MEM('o060514, 16'o000000);
`MEM('o060516, 16'o000000);
`MEM('o060520, 16'o000000);
`MEM('o060522, 16'o000000);
`MEM('o060524, 16'o000000);
`MEM('o060526, 16'o000000);
`MEM('o060530, 16'o000000);
`MEM('o060532, 16'o000000);
`MEM('o060534, 16'o000000);
`MEM('o060536, 16'o000000);
`MEM('o060540, 16'o000000);
`MEM('o060542, 16'o000000);
`MEM('o060544, 16'o000000);
`MEM('o060546, 16'o000000);
`MEM('o060550, 16'o000000);
`MEM('o060552, 16'o000000);
`MEM('o060554, 16'o000000);
`MEM('o060556, 16'o000000);
`MEM('o060560, 16'o000000);
`MEM('o060562, 16'o000000);
`MEM('o060564, 16'o000000);
`MEM('o060566, 16'o000000);
`MEM('o060570, 16'o000000);
`MEM('o060572, 16'o000000);
`MEM('o060574, 16'o000000);
`MEM('o060576, 16'o000000);
`MEM('o060600, 16'o000000);
`MEM('o060602, 16'o000000);
`MEM('o060604, 16'o000000);
`MEM('o060606, 16'o000000);
`MEM('o060610, 16'o000000);
`MEM('o060612, 16'o000000);
`MEM('o060614, 16'o000000);
`MEM('o060616, 16'o000000);
`MEM('o060620, 16'o000000);
`MEM('o060622, 16'o000000);
`MEM('o060624, 16'o000000);
`MEM('o060626, 16'o000000);
`MEM('o060630, 16'o000000);
`MEM('o060632, 16'o000000);
`MEM('o060634, 16'o000000);
`MEM('o060636, 16'o000000);
`MEM('o060640, 16'o000000);
`MEM('o060642, 16'o000000);
`MEM('o060644, 16'o000000);
`MEM('o060646, 16'o000000);
`MEM('o060650, 16'o000000);
`MEM('o060652, 16'o000000);
`MEM('o060654, 16'o000000);
`MEM('o060656, 16'o000000);
`MEM('o060660, 16'o000000);
`MEM('o060662, 16'o000000);
`MEM('o060664, 16'o000000);
`MEM('o060666, 16'o000000);
`MEM('o060670, 16'o000000);
`MEM('o060672, 16'o000000);
`MEM('o060674, 16'o000000);
`MEM('o060676, 16'o000000);
`MEM('o060700, 16'o000000);
`MEM('o060702, 16'o000000);
`MEM('o060704, 16'o000000);
`MEM('o060706, 16'o000000);
`MEM('o060710, 16'o000000);
`MEM('o060712, 16'o000000);
`MEM('o060714, 16'o000000);
`MEM('o060716, 16'o000000);
`MEM('o060720, 16'o000000);
`MEM('o060722, 16'o000000);
`MEM('o060724, 16'o000000);
`MEM('o060726, 16'o000000);
`MEM('o060730, 16'o000000);
`MEM('o060732, 16'o000000);
`MEM('o060734, 16'o000000);
`MEM('o060736, 16'o000000);
`MEM('o060740, 16'o000000);
`MEM('o060742, 16'o000000);
`MEM('o060744, 16'o000000);
`MEM('o060746, 16'o000000);
`MEM('o060750, 16'o000000);
`MEM('o060752, 16'o000000);
`MEM('o060754, 16'o000000);
`MEM('o060756, 16'o000000);
`MEM('o060760, 16'o000000);
`MEM('o060762, 16'o000000);
`MEM('o060764, 16'o000000);
`MEM('o060766, 16'o000000);
`MEM('o060770, 16'o000000);
`MEM('o060772, 16'o000000);
`MEM('o060774, 16'o000000);
`MEM('o060776, 16'o000000);
`MEM('o061000, 16'o000000);
`MEM('o061002, 16'o000000);
`MEM('o061004, 16'o000000);
`MEM('o061006, 16'o000000);
`MEM('o061010, 16'o000000);
`MEM('o061012, 16'o000000);
`MEM('o061014, 16'o000000);
`MEM('o061016, 16'o000000);
`MEM('o061020, 16'o000000);
`MEM('o061022, 16'o000000);
`MEM('o061024, 16'o000000);
`MEM('o061026, 16'o000000);
`MEM('o061030, 16'o000000);
`MEM('o061032, 16'o000000);
`MEM('o061034, 16'o000000);
`MEM('o061036, 16'o000000);
`MEM('o061040, 16'o000000);
`MEM('o061042, 16'o000000);
`MEM('o061044, 16'o000000);
`MEM('o061046, 16'o000000);
`MEM('o061050, 16'o000000);
`MEM('o061052, 16'o000000);
`MEM('o061054, 16'o000000);
`MEM('o061056, 16'o000000);
`MEM('o061060, 16'o000000);
`MEM('o061062, 16'o000000);
`MEM('o061064, 16'o000000);
`MEM('o061066, 16'o000000);
`MEM('o061070, 16'o000000);
`MEM('o061072, 16'o000000);
`MEM('o061074, 16'o000000);
`MEM('o061076, 16'o000000);
`MEM('o061100, 16'o000000);
`MEM('o061102, 16'o000000);
`MEM('o061104, 16'o000000);
`MEM('o061106, 16'o000000);
`MEM('o061110, 16'o000000);
`MEM('o061112, 16'o000000);
`MEM('o061114, 16'o000000);
`MEM('o061116, 16'o000000);
`MEM('o061120, 16'o000000);
`MEM('o061122, 16'o000000);
`MEM('o061124, 16'o000000);
`MEM('o061126, 16'o000000);
`MEM('o061130, 16'o000000);
`MEM('o061132, 16'o000000);
`MEM('o061134, 16'o000000);
`MEM('o061136, 16'o000000);
`MEM('o061140, 16'o000000);
`MEM('o061142, 16'o000000);
`MEM('o061144, 16'o000000);
`MEM('o061146, 16'o000000);
`MEM('o061150, 16'o000000);
`MEM('o061152, 16'o000000);
`MEM('o061154, 16'o000000);
`MEM('o061156, 16'o000000);
`MEM('o061160, 16'o000000);
`MEM('o061162, 16'o000000);
`MEM('o061164, 16'o000000);
`MEM('o061166, 16'o000000);
`MEM('o061170, 16'o000000);
`MEM('o061172, 16'o000000);
`MEM('o061174, 16'o000000);
`MEM('o061176, 16'o000000);
`MEM('o061200, 16'o000000);
`MEM('o061202, 16'o000000);
`MEM('o061204, 16'o000000);
`MEM('o061206, 16'o000000);
`MEM('o061210, 16'o000000);
`MEM('o061212, 16'o000000);
`MEM('o061214, 16'o000000);
`MEM('o061216, 16'o000000);
`MEM('o061220, 16'o000000);
`MEM('o061222, 16'o000000);
`MEM('o061224, 16'o000000);
`MEM('o061226, 16'o000000);
`MEM('o061230, 16'o000000);
`MEM('o061232, 16'o000000);
`MEM('o061234, 16'o000000);
`MEM('o061236, 16'o000000);
`MEM('o061240, 16'o000000);
`MEM('o061242, 16'o000000);
`MEM('o061244, 16'o000000);
`MEM('o061246, 16'o000000);
`MEM('o061250, 16'o000000);
`MEM('o061252, 16'o000000);
`MEM('o061254, 16'o000000);
`MEM('o061256, 16'o000000);
`MEM('o061260, 16'o000000);
`MEM('o061262, 16'o000000);
`MEM('o061264, 16'o000000);
`MEM('o061266, 16'o000000);
`MEM('o061270, 16'o000000);
`MEM('o061272, 16'o000000);
`MEM('o061274, 16'o000000);
`MEM('o061276, 16'o000000);
`MEM('o061300, 16'o000000);
`MEM('o061302, 16'o000000);
`MEM('o061304, 16'o000000);
`MEM('o061306, 16'o000000);
`MEM('o061310, 16'o000000);
`MEM('o061312, 16'o000000);
`MEM('o061314, 16'o000000);
`MEM('o061316, 16'o000000);
`MEM('o061320, 16'o000000);
`MEM('o061322, 16'o000000);
`MEM('o061324, 16'o000000);
`MEM('o061326, 16'o000000);
`MEM('o061330, 16'o000000);
`MEM('o061332, 16'o000000);
`MEM('o061334, 16'o000000);
`MEM('o061336, 16'o000000);
`MEM('o061340, 16'o000000);
`MEM('o061342, 16'o000000);
`MEM('o061344, 16'o000000);
`MEM('o061346, 16'o000000);
`MEM('o061350, 16'o000000);
`MEM('o061352, 16'o000000);
`MEM('o061354, 16'o000000);
`MEM('o061356, 16'o000000);
`MEM('o061360, 16'o000000);
`MEM('o061362, 16'o000000);
`MEM('o061364, 16'o000000);
`MEM('o061366, 16'o000000);
`MEM('o061370, 16'o000000);
`MEM('o061372, 16'o000000);
`MEM('o061374, 16'o000000);
`MEM('o061376, 16'o000000);
`MEM('o061400, 16'o000000);
`MEM('o061402, 16'o000000);
`MEM('o061404, 16'o000000);
`MEM('o061406, 16'o000000);
`MEM('o061410, 16'o000000);
`MEM('o061412, 16'o000000);
`MEM('o061414, 16'o000000);
`MEM('o061416, 16'o000000);
`MEM('o061420, 16'o000000);
`MEM('o061422, 16'o000000);
`MEM('o061424, 16'o000000);
`MEM('o061426, 16'o000000);
`MEM('o061430, 16'o000000);
`MEM('o061432, 16'o000000);
`MEM('o061434, 16'o000000);
`MEM('o061436, 16'o000000);
`MEM('o061440, 16'o000000);
`MEM('o061442, 16'o000000);
`MEM('o061444, 16'o000000);
`MEM('o061446, 16'o000000);
`MEM('o061450, 16'o000000);
`MEM('o061452, 16'o000000);
`MEM('o061454, 16'o000000);
`MEM('o061456, 16'o000000);
`MEM('o061460, 16'o000000);
`MEM('o061462, 16'o000000);
`MEM('o061464, 16'o000000);
`MEM('o061466, 16'o000000);
`MEM('o061470, 16'o000000);
`MEM('o061472, 16'o000000);
`MEM('o061474, 16'o000000);
`MEM('o061476, 16'o000000);
`MEM('o061500, 16'o000000);
`MEM('o061502, 16'o000000);
`MEM('o061504, 16'o000000);
`MEM('o061506, 16'o000000);
`MEM('o061510, 16'o000000);
`MEM('o061512, 16'o000000);
`MEM('o061514, 16'o000000);
`MEM('o061516, 16'o000000);
`MEM('o061520, 16'o000000);
`MEM('o061522, 16'o000000);
`MEM('o061524, 16'o000000);
`MEM('o061526, 16'o000000);
`MEM('o061530, 16'o000000);
`MEM('o061532, 16'o000000);
`MEM('o061534, 16'o000000);
`MEM('o061536, 16'o000000);
`MEM('o061540, 16'o000000);
`MEM('o061542, 16'o000000);
`MEM('o061544, 16'o000000);
`MEM('o061546, 16'o000000);
`MEM('o061550, 16'o000000);
`MEM('o061552, 16'o000000);
`MEM('o061554, 16'o000000);
`MEM('o061556, 16'o000000);
`MEM('o061560, 16'o000000);
`MEM('o061562, 16'o000000);
`MEM('o061564, 16'o000000);
`MEM('o061566, 16'o000000);
`MEM('o061570, 16'o000000);
`MEM('o061572, 16'o000000);
`MEM('o061574, 16'o000000);
`MEM('o061576, 16'o000000);
`MEM('o061600, 16'o000000);
`MEM('o061602, 16'o000000);
`MEM('o061604, 16'o000000);
`MEM('o061606, 16'o000000);
`MEM('o061610, 16'o000000);
`MEM('o061612, 16'o000000);
`MEM('o061614, 16'o000000);
`MEM('o061616, 16'o000000);
`MEM('o061620, 16'o000000);
`MEM('o061622, 16'o000000);
`MEM('o061624, 16'o000000);
`MEM('o061626, 16'o000000);
`MEM('o061630, 16'o000000);
`MEM('o061632, 16'o000000);
`MEM('o061634, 16'o000000);
`MEM('o061636, 16'o000000);
`MEM('o061640, 16'o000000);
`MEM('o061642, 16'o000000);
`MEM('o061644, 16'o000000);
`MEM('o061646, 16'o000000);
`MEM('o061650, 16'o000000);
`MEM('o061652, 16'o000000);
`MEM('o061654, 16'o000000);
`MEM('o061656, 16'o000000);
`MEM('o061660, 16'o000000);
`MEM('o061662, 16'o000000);
`MEM('o061664, 16'o000000);
`MEM('o061666, 16'o000000);
`MEM('o061670, 16'o000000);
`MEM('o061672, 16'o000000);
`MEM('o061674, 16'o000000);
`MEM('o061676, 16'o000000);
`MEM('o061700, 16'o000000);
`MEM('o061702, 16'o000000);
`MEM('o061704, 16'o000000);
`MEM('o061706, 16'o000000);
`MEM('o061710, 16'o000000);
`MEM('o061712, 16'o000000);
`MEM('o061714, 16'o000000);
`MEM('o061716, 16'o000000);
`MEM('o061720, 16'o000000);
`MEM('o061722, 16'o000000);
`MEM('o061724, 16'o000000);
`MEM('o061726, 16'o000000);
`MEM('o061730, 16'o000000);
`MEM('o061732, 16'o000000);
`MEM('o061734, 16'o000000);
`MEM('o061736, 16'o000000);
`MEM('o061740, 16'o000000);
`MEM('o061742, 16'o000000);
`MEM('o061744, 16'o000000);
`MEM('o061746, 16'o000000);
`MEM('o061750, 16'o000000);
`MEM('o061752, 16'o000000);
`MEM('o061754, 16'o000000);
`MEM('o061756, 16'o000000);
`MEM('o061760, 16'o000000);
`MEM('o061762, 16'o000000);
`MEM('o061764, 16'o000000);
`MEM('o061766, 16'o000000);
`MEM('o061770, 16'o000000);
`MEM('o061772, 16'o000000);
`MEM('o061774, 16'o000000);
`MEM('o061776, 16'o000000);
`MEM('o062000, 16'o000000);
`MEM('o062002, 16'o000000);
`MEM('o062004, 16'o000000);
`MEM('o062006, 16'o000000);
`MEM('o062010, 16'o000000);
`MEM('o062012, 16'o000000);
`MEM('o062014, 16'o000000);
`MEM('o062016, 16'o000000);
`MEM('o062020, 16'o000000);
`MEM('o062022, 16'o000000);
`MEM('o062024, 16'o000000);
`MEM('o062026, 16'o000000);
`MEM('o062030, 16'o000000);
`MEM('o062032, 16'o000000);
`MEM('o062034, 16'o000000);
`MEM('o062036, 16'o000000);
`MEM('o062040, 16'o000000);
`MEM('o062042, 16'o000000);
`MEM('o062044, 16'o000000);
`MEM('o062046, 16'o000000);
`MEM('o062050, 16'o000000);
`MEM('o062052, 16'o000000);
`MEM('o062054, 16'o000000);
`MEM('o062056, 16'o000000);
`MEM('o062060, 16'o000000);
`MEM('o062062, 16'o000000);
`MEM('o062064, 16'o000000);
`MEM('o062066, 16'o000000);
`MEM('o062070, 16'o000000);
`MEM('o062072, 16'o000000);
`MEM('o062074, 16'o000000);
`MEM('o062076, 16'o000000);
`MEM('o062100, 16'o000000);
`MEM('o062102, 16'o000000);
`MEM('o062104, 16'o000000);
`MEM('o062106, 16'o000000);
`MEM('o062110, 16'o000000);
`MEM('o062112, 16'o000000);
`MEM('o062114, 16'o000000);
`MEM('o062116, 16'o000000);
`MEM('o062120, 16'o000000);
`MEM('o062122, 16'o000000);
`MEM('o062124, 16'o000000);
`MEM('o062126, 16'o000000);
`MEM('o062130, 16'o000000);
`MEM('o062132, 16'o000000);
`MEM('o062134, 16'o000000);
`MEM('o062136, 16'o000000);
`MEM('o062140, 16'o000000);
`MEM('o062142, 16'o000000);
`MEM('o062144, 16'o000000);
`MEM('o062146, 16'o000000);
`MEM('o062150, 16'o000000);
`MEM('o062152, 16'o000000);
`MEM('o062154, 16'o000000);
`MEM('o062156, 16'o000000);
`MEM('o062160, 16'o000000);
`MEM('o062162, 16'o000000);
`MEM('o062164, 16'o000000);
`MEM('o062166, 16'o000000);
`MEM('o062170, 16'o000000);
`MEM('o062172, 16'o000000);
`MEM('o062174, 16'o000000);
`MEM('o062176, 16'o000000);
`MEM('o062200, 16'o000000);
`MEM('o062202, 16'o000000);
`MEM('o062204, 16'o000000);
`MEM('o062206, 16'o000000);
`MEM('o062210, 16'o000000);
`MEM('o062212, 16'o000000);
`MEM('o062214, 16'o000000);
`MEM('o062216, 16'o000000);
`MEM('o062220, 16'o000000);
`MEM('o062222, 16'o000000);
`MEM('o062224, 16'o000000);
`MEM('o062226, 16'o000000);
`MEM('o062230, 16'o000000);
`MEM('o062232, 16'o000000);
`MEM('o062234, 16'o000000);
`MEM('o062236, 16'o000000);
`MEM('o062240, 16'o000000);
`MEM('o062242, 16'o000000);
`MEM('o062244, 16'o000000);
`MEM('o062246, 16'o000000);
`MEM('o062250, 16'o000000);
`MEM('o062252, 16'o000000);
`MEM('o062254, 16'o000000);
`MEM('o062256, 16'o000000);
`MEM('o062260, 16'o000000);
`MEM('o062262, 16'o000000);
`MEM('o062264, 16'o000000);
`MEM('o062266, 16'o000000);
`MEM('o062270, 16'o000000);
`MEM('o062272, 16'o000000);
`MEM('o062274, 16'o000000);
`MEM('o062276, 16'o000000);
`MEM('o062300, 16'o000000);
`MEM('o062302, 16'o000000);
`MEM('o062304, 16'o000000);
`MEM('o062306, 16'o000000);
`MEM('o062310, 16'o000000);
`MEM('o062312, 16'o000000);
`MEM('o062314, 16'o000000);
`MEM('o062316, 16'o000000);
`MEM('o062320, 16'o000000);
`MEM('o062322, 16'o000000);
`MEM('o062324, 16'o000000);
`MEM('o062326, 16'o000000);
`MEM('o062330, 16'o000000);
`MEM('o062332, 16'o000000);
`MEM('o062334, 16'o000000);
`MEM('o062336, 16'o000000);
`MEM('o062340, 16'o000000);
`MEM('o062342, 16'o000000);
`MEM('o062344, 16'o000000);
`MEM('o062346, 16'o000000);
`MEM('o062350, 16'o000000);
`MEM('o062352, 16'o000000);
`MEM('o062354, 16'o000000);
`MEM('o062356, 16'o000000);
`MEM('o062360, 16'o000000);
`MEM('o062362, 16'o000000);
`MEM('o062364, 16'o000000);
`MEM('o062366, 16'o000000);
`MEM('o062370, 16'o000000);
`MEM('o062372, 16'o000000);
`MEM('o062374, 16'o000000);
`MEM('o062376, 16'o000000);
`MEM('o062400, 16'o000000);
`MEM('o062402, 16'o000000);
`MEM('o062404, 16'o000000);
`MEM('o062406, 16'o000000);
`MEM('o062410, 16'o000000);
`MEM('o062412, 16'o000000);
`MEM('o062414, 16'o000000);
`MEM('o062416, 16'o000000);
`MEM('o062420, 16'o000000);
`MEM('o062422, 16'o000000);
`MEM('o062424, 16'o000000);
`MEM('o062426, 16'o000000);
`MEM('o062430, 16'o000000);
`MEM('o062432, 16'o000000);
`MEM('o062434, 16'o000000);
`MEM('o062436, 16'o000000);
`MEM('o062440, 16'o000000);
`MEM('o062442, 16'o000000);
`MEM('o062444, 16'o000000);
`MEM('o062446, 16'o000000);
`MEM('o062450, 16'o000000);
`MEM('o062452, 16'o000000);
`MEM('o062454, 16'o000000);
`MEM('o062456, 16'o000000);
`MEM('o062460, 16'o000000);
`MEM('o062462, 16'o000000);
`MEM('o062464, 16'o000000);
`MEM('o062466, 16'o000000);
`MEM('o062470, 16'o000000);
`MEM('o062472, 16'o000000);
`MEM('o062474, 16'o000000);
`MEM('o062476, 16'o000000);
`MEM('o062500, 16'o000000);
`MEM('o062502, 16'o000000);
`MEM('o062504, 16'o000000);
`MEM('o062506, 16'o000000);
`MEM('o062510, 16'o000000);
`MEM('o062512, 16'o000000);
`MEM('o062514, 16'o000000);
`MEM('o062516, 16'o000000);
`MEM('o062520, 16'o000000);
`MEM('o062522, 16'o000000);
`MEM('o062524, 16'o000000);
`MEM('o062526, 16'o000000);
`MEM('o062530, 16'o000000);
`MEM('o062532, 16'o000000);
`MEM('o062534, 16'o000000);
`MEM('o062536, 16'o000000);
`MEM('o062540, 16'o000000);
`MEM('o062542, 16'o000000);
`MEM('o062544, 16'o000000);
`MEM('o062546, 16'o000000);
`MEM('o062550, 16'o000000);
`MEM('o062552, 16'o000000);
`MEM('o062554, 16'o000000);
`MEM('o062556, 16'o000000);
`MEM('o062560, 16'o000000);
`MEM('o062562, 16'o000000);
`MEM('o062564, 16'o000000);
`MEM('o062566, 16'o000000);
`MEM('o062570, 16'o000000);
`MEM('o062572, 16'o000000);
`MEM('o062574, 16'o000000);
`MEM('o062576, 16'o000000);
`MEM('o062600, 16'o000000);
`MEM('o062602, 16'o000000);
`MEM('o062604, 16'o000000);
`MEM('o062606, 16'o000000);
`MEM('o062610, 16'o000000);
`MEM('o062612, 16'o000000);
`MEM('o062614, 16'o000000);
`MEM('o062616, 16'o000000);
`MEM('o062620, 16'o000000);
`MEM('o062622, 16'o000000);
`MEM('o062624, 16'o000000);
`MEM('o062626, 16'o000000);
`MEM('o062630, 16'o000000);
`MEM('o062632, 16'o000000);
`MEM('o062634, 16'o000000);
`MEM('o062636, 16'o000000);
`MEM('o062640, 16'o000000);
`MEM('o062642, 16'o000000);
`MEM('o062644, 16'o000000);
`MEM('o062646, 16'o000000);
`MEM('o062650, 16'o000000);
`MEM('o062652, 16'o000000);
`MEM('o062654, 16'o000000);
`MEM('o062656, 16'o000000);
`MEM('o062660, 16'o000000);
`MEM('o062662, 16'o000000);
`MEM('o062664, 16'o000000);
`MEM('o062666, 16'o000000);
`MEM('o062670, 16'o000000);
`MEM('o062672, 16'o000000);
`MEM('o062674, 16'o000000);
`MEM('o062676, 16'o000000);
`MEM('o062700, 16'o000000);
`MEM('o062702, 16'o000000);
`MEM('o062704, 16'o000000);
`MEM('o062706, 16'o000000);
`MEM('o062710, 16'o000000);
`MEM('o062712, 16'o000000);
`MEM('o062714, 16'o000000);
`MEM('o062716, 16'o000000);
`MEM('o062720, 16'o000000);
`MEM('o062722, 16'o000000);
`MEM('o062724, 16'o000000);
`MEM('o062726, 16'o000000);
`MEM('o062730, 16'o000000);
`MEM('o062732, 16'o000000);
`MEM('o062734, 16'o000000);
`MEM('o062736, 16'o000000);
`MEM('o062740, 16'o000000);
`MEM('o062742, 16'o000000);
`MEM('o062744, 16'o000000);
`MEM('o062746, 16'o000000);
`MEM('o062750, 16'o000000);
`MEM('o062752, 16'o000000);
`MEM('o062754, 16'o000000);
`MEM('o062756, 16'o000000);
`MEM('o062760, 16'o000000);
`MEM('o062762, 16'o000000);
`MEM('o062764, 16'o000000);
`MEM('o062766, 16'o000000);
`MEM('o062770, 16'o000000);
`MEM('o062772, 16'o000000);
`MEM('o062774, 16'o000000);
`MEM('o062776, 16'o000000);
`MEM('o063000, 16'o000000);
`MEM('o063002, 16'o000000);
`MEM('o063004, 16'o000000);
`MEM('o063006, 16'o000000);
`MEM('o063010, 16'o000000);
`MEM('o063012, 16'o000000);
`MEM('o063014, 16'o000000);
`MEM('o063016, 16'o000000);
`MEM('o063020, 16'o000000);
`MEM('o063022, 16'o000000);
`MEM('o063024, 16'o000000);
`MEM('o063026, 16'o000000);
`MEM('o063030, 16'o000000);
`MEM('o063032, 16'o000000);
`MEM('o063034, 16'o000000);
`MEM('o063036, 16'o000000);
`MEM('o063040, 16'o000000);
`MEM('o063042, 16'o000000);
`MEM('o063044, 16'o000000);
`MEM('o063046, 16'o000000);
`MEM('o063050, 16'o000000);
`MEM('o063052, 16'o000000);
`MEM('o063054, 16'o000000);
`MEM('o063056, 16'o000000);
`MEM('o063060, 16'o000000);
`MEM('o063062, 16'o000000);
`MEM('o063064, 16'o000000);
`MEM('o063066, 16'o000000);
`MEM('o063070, 16'o000000);
`MEM('o063072, 16'o000000);
`MEM('o063074, 16'o000000);
`MEM('o063076, 16'o000000);
`MEM('o063100, 16'o000000);
`MEM('o063102, 16'o000000);
`MEM('o063104, 16'o000000);
`MEM('o063106, 16'o000000);
`MEM('o063110, 16'o000000);
`MEM('o063112, 16'o000000);
`MEM('o063114, 16'o000000);
`MEM('o063116, 16'o000000);
`MEM('o063120, 16'o000000);
`MEM('o063122, 16'o000000);
`MEM('o063124, 16'o000000);
`MEM('o063126, 16'o000000);
`MEM('o063130, 16'o000000);
`MEM('o063132, 16'o000000);
`MEM('o063134, 16'o000000);
`MEM('o063136, 16'o000000);
`MEM('o063140, 16'o000000);
`MEM('o063142, 16'o000000);
`MEM('o063144, 16'o000000);
`MEM('o063146, 16'o000000);
`MEM('o063150, 16'o000000);
`MEM('o063152, 16'o000000);
`MEM('o063154, 16'o000000);
`MEM('o063156, 16'o000000);
`MEM('o063160, 16'o000000);
`MEM('o063162, 16'o000000);
`MEM('o063164, 16'o000000);
`MEM('o063166, 16'o000000);
`MEM('o063170, 16'o000000);
`MEM('o063172, 16'o000000);
`MEM('o063174, 16'o000000);
`MEM('o063176, 16'o000000);
`MEM('o063200, 16'o000000);
`MEM('o063202, 16'o000000);
`MEM('o063204, 16'o000000);
`MEM('o063206, 16'o000000);
`MEM('o063210, 16'o000000);
`MEM('o063212, 16'o000000);
`MEM('o063214, 16'o000000);
`MEM('o063216, 16'o000000);
`MEM('o063220, 16'o000000);
`MEM('o063222, 16'o000000);
`MEM('o063224, 16'o000000);
`MEM('o063226, 16'o000000);
`MEM('o063230, 16'o000000);
`MEM('o063232, 16'o000000);
`MEM('o063234, 16'o000000);
`MEM('o063236, 16'o000000);
`MEM('o063240, 16'o000000);
`MEM('o063242, 16'o000000);
`MEM('o063244, 16'o000000);
`MEM('o063246, 16'o000000);
`MEM('o063250, 16'o000000);
`MEM('o063252, 16'o000000);
`MEM('o063254, 16'o000000);
`MEM('o063256, 16'o000000);
`MEM('o063260, 16'o000000);
`MEM('o063262, 16'o000000);
`MEM('o063264, 16'o000000);
`MEM('o063266, 16'o000000);
`MEM('o063270, 16'o000000);
`MEM('o063272, 16'o000000);
`MEM('o063274, 16'o000000);
`MEM('o063276, 16'o000000);
`MEM('o063300, 16'o000000);
`MEM('o063302, 16'o000000);
`MEM('o063304, 16'o000000);
`MEM('o063306, 16'o000000);
`MEM('o063310, 16'o000000);
`MEM('o063312, 16'o000000);
`MEM('o063314, 16'o000000);
`MEM('o063316, 16'o000000);
`MEM('o063320, 16'o000000);
`MEM('o063322, 16'o000000);
`MEM('o063324, 16'o000000);
`MEM('o063326, 16'o000000);
`MEM('o063330, 16'o000000);
`MEM('o063332, 16'o000000);
`MEM('o063334, 16'o000000);
`MEM('o063336, 16'o000000);
`MEM('o063340, 16'o000000);
`MEM('o063342, 16'o000000);
`MEM('o063344, 16'o000000);
`MEM('o063346, 16'o000000);
`MEM('o063350, 16'o000000);
`MEM('o063352, 16'o000000);
`MEM('o063354, 16'o000000);
`MEM('o063356, 16'o000000);
`MEM('o063360, 16'o000000);
`MEM('o063362, 16'o000000);
`MEM('o063364, 16'o000000);
`MEM('o063366, 16'o000000);
`MEM('o063370, 16'o000000);
`MEM('o063372, 16'o000000);
`MEM('o063374, 16'o000000);
`MEM('o063376, 16'o000000);
`MEM('o063400, 16'o000000);
`MEM('o063402, 16'o000000);
`MEM('o063404, 16'o000000);
`MEM('o063406, 16'o000000);
`MEM('o063410, 16'o000000);
`MEM('o063412, 16'o000000);
`MEM('o063414, 16'o000000);
`MEM('o063416, 16'o000000);
`MEM('o063420, 16'o000000);
`MEM('o063422, 16'o000000);
`MEM('o063424, 16'o000000);
`MEM('o063426, 16'o000000);
`MEM('o063430, 16'o000000);
`MEM('o063432, 16'o000000);
`MEM('o063434, 16'o000000);
`MEM('o063436, 16'o000000);
`MEM('o063440, 16'o000000);
`MEM('o063442, 16'o000000);
`MEM('o063444, 16'o000000);
`MEM('o063446, 16'o000000);
`MEM('o063450, 16'o000000);
`MEM('o063452, 16'o000000);
`MEM('o063454, 16'o000000);
`MEM('o063456, 16'o000000);
`MEM('o063460, 16'o000000);
`MEM('o063462, 16'o000000);
`MEM('o063464, 16'o000000);
`MEM('o063466, 16'o000000);
`MEM('o063470, 16'o000000);
`MEM('o063472, 16'o000000);
`MEM('o063474, 16'o000000);
`MEM('o063476, 16'o000000);
`MEM('o063500, 16'o000000);
`MEM('o063502, 16'o000000);
`MEM('o063504, 16'o000000);
`MEM('o063506, 16'o000000);
`MEM('o063510, 16'o000000);
`MEM('o063512, 16'o000000);
`MEM('o063514, 16'o000000);
`MEM('o063516, 16'o000000);
`MEM('o063520, 16'o000000);
`MEM('o063522, 16'o000000);
`MEM('o063524, 16'o000000);
`MEM('o063526, 16'o000000);
`MEM('o063530, 16'o000000);
`MEM('o063532, 16'o000000);
`MEM('o063534, 16'o000000);
`MEM('o063536, 16'o000000);
`MEM('o063540, 16'o000000);
`MEM('o063542, 16'o000000);
`MEM('o063544, 16'o000000);
`MEM('o063546, 16'o000000);
`MEM('o063550, 16'o000000);
`MEM('o063552, 16'o000000);
`MEM('o063554, 16'o000000);
`MEM('o063556, 16'o000000);
`MEM('o063560, 16'o000000);
`MEM('o063562, 16'o000000);
`MEM('o063564, 16'o000000);
`MEM('o063566, 16'o000000);
`MEM('o063570, 16'o000000);
`MEM('o063572, 16'o000000);
`MEM('o063574, 16'o000000);
`MEM('o063576, 16'o000000);
`MEM('o063600, 16'o000000);
`MEM('o063602, 16'o000000);
`MEM('o063604, 16'o000000);
`MEM('o063606, 16'o000000);
`MEM('o063610, 16'o000000);
`MEM('o063612, 16'o000000);
`MEM('o063614, 16'o000000);
`MEM('o063616, 16'o000000);
`MEM('o063620, 16'o000000);
`MEM('o063622, 16'o000000);
`MEM('o063624, 16'o000000);
`MEM('o063626, 16'o000000);
`MEM('o063630, 16'o000000);
`MEM('o063632, 16'o000000);
`MEM('o063634, 16'o000000);
`MEM('o063636, 16'o000000);
`MEM('o063640, 16'o000000);
`MEM('o063642, 16'o000000);
`MEM('o063644, 16'o000000);
`MEM('o063646, 16'o000000);
`MEM('o063650, 16'o000000);
`MEM('o063652, 16'o000000);
`MEM('o063654, 16'o000000);
`MEM('o063656, 16'o000000);
`MEM('o063660, 16'o000000);
`MEM('o063662, 16'o000000);
`MEM('o063664, 16'o000000);
`MEM('o063666, 16'o000000);
`MEM('o063670, 16'o000000);
`MEM('o063672, 16'o000000);
`MEM('o063674, 16'o000000);
`MEM('o063676, 16'o000000);
`MEM('o063700, 16'o000000);
`MEM('o063702, 16'o000000);
`MEM('o063704, 16'o000000);
`MEM('o063706, 16'o000000);
`MEM('o063710, 16'o000000);
`MEM('o063712, 16'o000000);
`MEM('o063714, 16'o000000);
`MEM('o063716, 16'o000000);
`MEM('o063720, 16'o000000);
`MEM('o063722, 16'o000000);
`MEM('o063724, 16'o000000);
`MEM('o063726, 16'o000000);
`MEM('o063730, 16'o000000);
`MEM('o063732, 16'o000000);
`MEM('o063734, 16'o000000);
`MEM('o063736, 16'o000000);
`MEM('o063740, 16'o000000);
`MEM('o063742, 16'o000000);
`MEM('o063744, 16'o000000);
`MEM('o063746, 16'o000000);
`MEM('o063750, 16'o000000);
`MEM('o063752, 16'o000000);
`MEM('o063754, 16'o000000);
`MEM('o063756, 16'o000000);
`MEM('o063760, 16'o000000);
`MEM('o063762, 16'o000000);
`MEM('o063764, 16'o000000);
`MEM('o063766, 16'o000000);
`MEM('o063770, 16'o000000);
`MEM('o063772, 16'o000000);
`MEM('o063774, 16'o000000);
`MEM('o063776, 16'o000000);
`MEM('o064000, 16'o000000);
`MEM('o064002, 16'o000000);
`MEM('o064004, 16'o000000);
`MEM('o064006, 16'o000000);
`MEM('o064010, 16'o000000);
`MEM('o064012, 16'o000000);
`MEM('o064014, 16'o000000);
`MEM('o064016, 16'o000000);
`MEM('o064020, 16'o000000);
`MEM('o064022, 16'o000000);
`MEM('o064024, 16'o000000);
`MEM('o064026, 16'o000000);
`MEM('o064030, 16'o000000);
`MEM('o064032, 16'o000000);
`MEM('o064034, 16'o000000);
`MEM('o064036, 16'o000000);
`MEM('o064040, 16'o000000);
`MEM('o064042, 16'o000000);
`MEM('o064044, 16'o000000);
`MEM('o064046, 16'o000000);
`MEM('o064050, 16'o000000);
`MEM('o064052, 16'o000000);
`MEM('o064054, 16'o000000);
`MEM('o064056, 16'o000000);
`MEM('o064060, 16'o000000);
`MEM('o064062, 16'o000000);
`MEM('o064064, 16'o000000);
`MEM('o064066, 16'o000000);
`MEM('o064070, 16'o000000);
`MEM('o064072, 16'o000000);
`MEM('o064074, 16'o000000);
`MEM('o064076, 16'o000000);
`MEM('o064100, 16'o000000);
`MEM('o064102, 16'o000000);
`MEM('o064104, 16'o000000);
`MEM('o064106, 16'o000000);
`MEM('o064110, 16'o000000);
`MEM('o064112, 16'o000000);
`MEM('o064114, 16'o000000);
`MEM('o064116, 16'o000000);
`MEM('o064120, 16'o000000);
`MEM('o064122, 16'o000000);
`MEM('o064124, 16'o000000);
`MEM('o064126, 16'o000000);
`MEM('o064130, 16'o000000);
`MEM('o064132, 16'o000000);
`MEM('o064134, 16'o000000);
`MEM('o064136, 16'o000000);
`MEM('o064140, 16'o000000);
`MEM('o064142, 16'o000000);
`MEM('o064144, 16'o000000);
`MEM('o064146, 16'o000000);
`MEM('o064150, 16'o000000);
`MEM('o064152, 16'o000000);
`MEM('o064154, 16'o000000);
`MEM('o064156, 16'o000000);
`MEM('o064160, 16'o000000);
`MEM('o064162, 16'o000000);
`MEM('o064164, 16'o000000);
`MEM('o064166, 16'o000000);
`MEM('o064170, 16'o000000);
`MEM('o064172, 16'o000000);
`MEM('o064174, 16'o000000);
`MEM('o064176, 16'o000000);
`MEM('o064200, 16'o000000);
`MEM('o064202, 16'o000000);
`MEM('o064204, 16'o000000);
`MEM('o064206, 16'o000000);
`MEM('o064210, 16'o000000);
`MEM('o064212, 16'o000000);
`MEM('o064214, 16'o000000);
`MEM('o064216, 16'o000000);
`MEM('o064220, 16'o000000);
`MEM('o064222, 16'o000000);
`MEM('o064224, 16'o000000);
`MEM('o064226, 16'o000000);
`MEM('o064230, 16'o000000);
`MEM('o064232, 16'o000000);
`MEM('o064234, 16'o000000);
`MEM('o064236, 16'o000000);
`MEM('o064240, 16'o000000);
`MEM('o064242, 16'o000000);
`MEM('o064244, 16'o000000);
`MEM('o064246, 16'o000000);
`MEM('o064250, 16'o000000);
`MEM('o064252, 16'o000000);
`MEM('o064254, 16'o000000);
`MEM('o064256, 16'o000000);
`MEM('o064260, 16'o000000);
`MEM('o064262, 16'o000000);
`MEM('o064264, 16'o000000);
`MEM('o064266, 16'o000000);
`MEM('o064270, 16'o000000);
`MEM('o064272, 16'o000000);
`MEM('o064274, 16'o000000);
`MEM('o064276, 16'o000000);
`MEM('o064300, 16'o000000);
`MEM('o064302, 16'o000000);
`MEM('o064304, 16'o000000);
`MEM('o064306, 16'o000000);
`MEM('o064310, 16'o000000);
`MEM('o064312, 16'o000000);
`MEM('o064314, 16'o000000);
`MEM('o064316, 16'o000000);
`MEM('o064320, 16'o000000);
`MEM('o064322, 16'o000000);
`MEM('o064324, 16'o000000);
`MEM('o064326, 16'o000000);
`MEM('o064330, 16'o000000);
`MEM('o064332, 16'o000000);
`MEM('o064334, 16'o000000);
`MEM('o064336, 16'o000000);
`MEM('o064340, 16'o000000);
`MEM('o064342, 16'o000000);
`MEM('o064344, 16'o000000);
`MEM('o064346, 16'o000000);
`MEM('o064350, 16'o000000);
`MEM('o064352, 16'o000000);
`MEM('o064354, 16'o000000);
`MEM('o064356, 16'o000000);
`MEM('o064360, 16'o000000);
`MEM('o064362, 16'o000000);
`MEM('o064364, 16'o000000);
`MEM('o064366, 16'o000000);
`MEM('o064370, 16'o000000);
`MEM('o064372, 16'o000000);
`MEM('o064374, 16'o000000);
`MEM('o064376, 16'o000000);
`MEM('o064400, 16'o000000);
`MEM('o064402, 16'o000000);
`MEM('o064404, 16'o000000);
`MEM('o064406, 16'o000000);
`MEM('o064410, 16'o000000);
`MEM('o064412, 16'o000000);
`MEM('o064414, 16'o000000);
`MEM('o064416, 16'o000000);
`MEM('o064420, 16'o000000);
`MEM('o064422, 16'o000000);
`MEM('o064424, 16'o000000);
`MEM('o064426, 16'o000000);
`MEM('o064430, 16'o000000);
`MEM('o064432, 16'o000000);
`MEM('o064434, 16'o000000);
`MEM('o064436, 16'o000000);
`MEM('o064440, 16'o000000);
`MEM('o064442, 16'o000000);
`MEM('o064444, 16'o000000);
`MEM('o064446, 16'o000000);
`MEM('o064450, 16'o000000);
`MEM('o064452, 16'o000000);
`MEM('o064454, 16'o000000);
`MEM('o064456, 16'o000000);
`MEM('o064460, 16'o000000);
`MEM('o064462, 16'o000000);
`MEM('o064464, 16'o000000);
`MEM('o064466, 16'o000000);
`MEM('o064470, 16'o000000);
`MEM('o064472, 16'o000000);
`MEM('o064474, 16'o000000);
`MEM('o064476, 16'o000000);
`MEM('o064500, 16'o000000);
`MEM('o064502, 16'o000000);
`MEM('o064504, 16'o000000);
`MEM('o064506, 16'o000000);
`MEM('o064510, 16'o000000);
`MEM('o064512, 16'o000000);
`MEM('o064514, 16'o000000);
`MEM('o064516, 16'o000000);
`MEM('o064520, 16'o000000);
`MEM('o064522, 16'o000000);
`MEM('o064524, 16'o000000);
`MEM('o064526, 16'o000000);
`MEM('o064530, 16'o000000);
`MEM('o064532, 16'o000000);
`MEM('o064534, 16'o000000);
`MEM('o064536, 16'o000000);
`MEM('o064540, 16'o000000);
`MEM('o064542, 16'o000000);
`MEM('o064544, 16'o000000);
`MEM('o064546, 16'o000000);
`MEM('o064550, 16'o000000);
`MEM('o064552, 16'o000000);
`MEM('o064554, 16'o000000);
`MEM('o064556, 16'o000000);
`MEM('o064560, 16'o000000);
`MEM('o064562, 16'o000000);
`MEM('o064564, 16'o000000);
`MEM('o064566, 16'o000000);
`MEM('o064570, 16'o000000);
`MEM('o064572, 16'o000000);
`MEM('o064574, 16'o000000);
`MEM('o064576, 16'o000000);
`MEM('o064600, 16'o000000);
`MEM('o064602, 16'o000000);
`MEM('o064604, 16'o000000);
`MEM('o064606, 16'o000000);
`MEM('o064610, 16'o000000);
`MEM('o064612, 16'o000000);
`MEM('o064614, 16'o000000);
`MEM('o064616, 16'o000000);
`MEM('o064620, 16'o000000);
`MEM('o064622, 16'o000000);
`MEM('o064624, 16'o000000);
`MEM('o064626, 16'o000000);
`MEM('o064630, 16'o000000);
`MEM('o064632, 16'o000000);
`MEM('o064634, 16'o000000);
`MEM('o064636, 16'o000000);
`MEM('o064640, 16'o000000);
`MEM('o064642, 16'o000000);
`MEM('o064644, 16'o000000);
`MEM('o064646, 16'o000000);
`MEM('o064650, 16'o000000);
`MEM('o064652, 16'o000000);
`MEM('o064654, 16'o000000);
`MEM('o064656, 16'o000000);
`MEM('o064660, 16'o000000);
`MEM('o064662, 16'o000000);
`MEM('o064664, 16'o000000);
`MEM('o064666, 16'o000000);
`MEM('o064670, 16'o000000);
`MEM('o064672, 16'o000000);
`MEM('o064674, 16'o000000);
`MEM('o064676, 16'o000000);
`MEM('o064700, 16'o000000);
`MEM('o064702, 16'o000000);
`MEM('o064704, 16'o000000);
`MEM('o064706, 16'o000000);
`MEM('o064710, 16'o000000);
`MEM('o064712, 16'o000000);
`MEM('o064714, 16'o000000);
`MEM('o064716, 16'o000000);
`MEM('o064720, 16'o000000);
`MEM('o064722, 16'o000000);
`MEM('o064724, 16'o000000);
`MEM('o064726, 16'o000000);
`MEM('o064730, 16'o000000);
`MEM('o064732, 16'o000000);
`MEM('o064734, 16'o000000);
`MEM('o064736, 16'o000000);
`MEM('o064740, 16'o000000);
`MEM('o064742, 16'o000000);
`MEM('o064744, 16'o000000);
`MEM('o064746, 16'o000000);
`MEM('o064750, 16'o000000);
`MEM('o064752, 16'o000000);
`MEM('o064754, 16'o000000);
`MEM('o064756, 16'o000000);
`MEM('o064760, 16'o000000);
`MEM('o064762, 16'o000000);
`MEM('o064764, 16'o000000);
`MEM('o064766, 16'o000000);
`MEM('o064770, 16'o000000);
`MEM('o064772, 16'o000000);
`MEM('o064774, 16'o000000);
`MEM('o064776, 16'o000000);
`MEM('o065000, 16'o000000);
`MEM('o065002, 16'o000000);
`MEM('o065004, 16'o000000);
`MEM('o065006, 16'o000000);
`MEM('o065010, 16'o000000);
`MEM('o065012, 16'o000000);
`MEM('o065014, 16'o000000);
`MEM('o065016, 16'o000000);
`MEM('o065020, 16'o000000);
`MEM('o065022, 16'o000000);
`MEM('o065024, 16'o000000);
`MEM('o065026, 16'o000000);
`MEM('o065030, 16'o000000);
`MEM('o065032, 16'o000000);
`MEM('o065034, 16'o000000);
`MEM('o065036, 16'o000000);
`MEM('o065040, 16'o000000);
`MEM('o065042, 16'o000000);
`MEM('o065044, 16'o000000);
`MEM('o065046, 16'o000000);
`MEM('o065050, 16'o000000);
`MEM('o065052, 16'o000000);
`MEM('o065054, 16'o000000);
`MEM('o065056, 16'o000000);
`MEM('o065060, 16'o000000);
`MEM('o065062, 16'o000000);
`MEM('o065064, 16'o000000);
`MEM('o065066, 16'o000000);
`MEM('o065070, 16'o000000);
`MEM('o065072, 16'o000000);
`MEM('o065074, 16'o000000);
`MEM('o065076, 16'o000000);
`MEM('o065100, 16'o000000);
`MEM('o065102, 16'o000000);
`MEM('o065104, 16'o000000);
`MEM('o065106, 16'o000000);
`MEM('o065110, 16'o000000);
`MEM('o065112, 16'o000000);
`MEM('o065114, 16'o000000);
`MEM('o065116, 16'o000000);
`MEM('o065120, 16'o000000);
`MEM('o065122, 16'o000000);
`MEM('o065124, 16'o000000);
`MEM('o065126, 16'o000000);
`MEM('o065130, 16'o000000);
`MEM('o065132, 16'o000000);
`MEM('o065134, 16'o000000);
`MEM('o065136, 16'o000000);
`MEM('o065140, 16'o000000);
`MEM('o065142, 16'o000000);
`MEM('o065144, 16'o000000);
`MEM('o065146, 16'o000000);
`MEM('o065150, 16'o000000);
`MEM('o065152, 16'o000000);
`MEM('o065154, 16'o000000);
`MEM('o065156, 16'o000000);
`MEM('o065160, 16'o000000);
`MEM('o065162, 16'o000000);
`MEM('o065164, 16'o000000);
`MEM('o065166, 16'o000000);
`MEM('o065170, 16'o000000);
`MEM('o065172, 16'o000000);
`MEM('o065174, 16'o000000);
`MEM('o065176, 16'o000000);
`MEM('o065200, 16'o000000);
`MEM('o065202, 16'o000000);
`MEM('o065204, 16'o000000);
`MEM('o065206, 16'o000000);
`MEM('o065210, 16'o000000);
`MEM('o065212, 16'o000000);
`MEM('o065214, 16'o000000);
`MEM('o065216, 16'o000000);
`MEM('o065220, 16'o000000);
`MEM('o065222, 16'o000000);
`MEM('o065224, 16'o000000);
`MEM('o065226, 16'o000000);
`MEM('o065230, 16'o000000);
`MEM('o065232, 16'o000000);
`MEM('o065234, 16'o000000);
`MEM('o065236, 16'o000000);
`MEM('o065240, 16'o000000);
`MEM('o065242, 16'o000000);
`MEM('o065244, 16'o000000);
`MEM('o065246, 16'o000000);
`MEM('o065250, 16'o000000);
`MEM('o065252, 16'o000000);
`MEM('o065254, 16'o000000);
`MEM('o065256, 16'o000000);
`MEM('o065260, 16'o000000);
`MEM('o065262, 16'o000000);
`MEM('o065264, 16'o000000);
`MEM('o065266, 16'o000000);
`MEM('o065270, 16'o000000);
`MEM('o065272, 16'o000000);
`MEM('o065274, 16'o000000);
`MEM('o065276, 16'o000000);
`MEM('o065300, 16'o000000);
`MEM('o065302, 16'o000000);
`MEM('o065304, 16'o000000);
`MEM('o065306, 16'o000000);
`MEM('o065310, 16'o000000);
`MEM('o065312, 16'o000000);
`MEM('o065314, 16'o000000);
`MEM('o065316, 16'o000000);
`MEM('o065320, 16'o000000);
`MEM('o065322, 16'o000000);
`MEM('o065324, 16'o000000);
`MEM('o065326, 16'o000000);
`MEM('o065330, 16'o000000);
`MEM('o065332, 16'o000000);
`MEM('o065334, 16'o000000);
`MEM('o065336, 16'o000000);
`MEM('o065340, 16'o000000);
`MEM('o065342, 16'o000000);
`MEM('o065344, 16'o000000);
`MEM('o065346, 16'o000000);
`MEM('o065350, 16'o000000);
`MEM('o065352, 16'o000000);
`MEM('o065354, 16'o000000);
`MEM('o065356, 16'o000000);
`MEM('o065360, 16'o000000);
`MEM('o065362, 16'o000000);
`MEM('o065364, 16'o000000);
`MEM('o065366, 16'o000000);
`MEM('o065370, 16'o000000);
`MEM('o065372, 16'o000000);
`MEM('o065374, 16'o000000);
`MEM('o065376, 16'o000000);
`MEM('o065400, 16'o000000);
`MEM('o065402, 16'o000000);
`MEM('o065404, 16'o000000);
`MEM('o065406, 16'o000000);
`MEM('o065410, 16'o000000);
`MEM('o065412, 16'o000000);
`MEM('o065414, 16'o000000);
`MEM('o065416, 16'o000000);
`MEM('o065420, 16'o000000);
`MEM('o065422, 16'o000000);
`MEM('o065424, 16'o000000);
`MEM('o065426, 16'o000000);
`MEM('o065430, 16'o000000);
`MEM('o065432, 16'o000000);
`MEM('o065434, 16'o000000);
`MEM('o065436, 16'o000000);
`MEM('o065440, 16'o000000);
`MEM('o065442, 16'o000000);
`MEM('o065444, 16'o000000);
`MEM('o065446, 16'o000000);
`MEM('o065450, 16'o000000);
`MEM('o065452, 16'o000000);
`MEM('o065454, 16'o000000);
`MEM('o065456, 16'o000000);
`MEM('o065460, 16'o000000);
`MEM('o065462, 16'o000000);
`MEM('o065464, 16'o000000);
`MEM('o065466, 16'o000000);
`MEM('o065470, 16'o000000);
`MEM('o065472, 16'o000000);
`MEM('o065474, 16'o000000);
`MEM('o065476, 16'o000000);
`MEM('o065500, 16'o000000);
`MEM('o065502, 16'o000000);
`MEM('o065504, 16'o000000);
`MEM('o065506, 16'o000000);
`MEM('o065510, 16'o000000);
`MEM('o065512, 16'o000000);
`MEM('o065514, 16'o000000);
`MEM('o065516, 16'o000000);
`MEM('o065520, 16'o000000);
`MEM('o065522, 16'o000000);
`MEM('o065524, 16'o000000);
`MEM('o065526, 16'o000000);
`MEM('o065530, 16'o000000);
`MEM('o065532, 16'o000000);
`MEM('o065534, 16'o000000);
`MEM('o065536, 16'o000000);
`MEM('o065540, 16'o000000);
`MEM('o065542, 16'o000000);
`MEM('o065544, 16'o000000);
`MEM('o065546, 16'o000000);
`MEM('o065550, 16'o000000);
`MEM('o065552, 16'o000000);
`MEM('o065554, 16'o000000);
`MEM('o065556, 16'o000000);
`MEM('o065560, 16'o000000);
`MEM('o065562, 16'o000000);
`MEM('o065564, 16'o000000);
`MEM('o065566, 16'o000000);
`MEM('o065570, 16'o000000);
`MEM('o065572, 16'o000000);
`MEM('o065574, 16'o000000);
`MEM('o065576, 16'o000000);
`MEM('o065600, 16'o000000);
`MEM('o065602, 16'o000000);
`MEM('o065604, 16'o000000);
`MEM('o065606, 16'o000000);
`MEM('o065610, 16'o000000);
`MEM('o065612, 16'o000000);
`MEM('o065614, 16'o000000);
`MEM('o065616, 16'o000000);
`MEM('o065620, 16'o000000);
`MEM('o065622, 16'o000000);
`MEM('o065624, 16'o000000);
`MEM('o065626, 16'o000000);
`MEM('o065630, 16'o000000);
`MEM('o065632, 16'o000000);
`MEM('o065634, 16'o000000);
`MEM('o065636, 16'o000000);
`MEM('o065640, 16'o000000);
`MEM('o065642, 16'o000000);
`MEM('o065644, 16'o000000);
`MEM('o065646, 16'o000000);
`MEM('o065650, 16'o000000);
`MEM('o065652, 16'o000000);
`MEM('o065654, 16'o000000);
`MEM('o065656, 16'o000000);
`MEM('o065660, 16'o000000);
`MEM('o065662, 16'o000000);
`MEM('o065664, 16'o000000);
`MEM('o065666, 16'o000000);
`MEM('o065670, 16'o000000);
`MEM('o065672, 16'o000000);
`MEM('o065674, 16'o000000);
`MEM('o065676, 16'o000000);
`MEM('o065700, 16'o000000);
`MEM('o065702, 16'o000000);
`MEM('o065704, 16'o000000);
`MEM('o065706, 16'o000000);
`MEM('o065710, 16'o000000);
`MEM('o065712, 16'o000000);
`MEM('o065714, 16'o000000);
`MEM('o065716, 16'o000000);
`MEM('o065720, 16'o000000);
`MEM('o065722, 16'o000000);
`MEM('o065724, 16'o000000);
`MEM('o065726, 16'o000000);
`MEM('o065730, 16'o000000);
`MEM('o065732, 16'o000000);
`MEM('o065734, 16'o000000);
`MEM('o065736, 16'o000000);
`MEM('o065740, 16'o000000);
`MEM('o065742, 16'o000000);
`MEM('o065744, 16'o000000);
`MEM('o065746, 16'o000000);
`MEM('o065750, 16'o000000);
`MEM('o065752, 16'o000000);
`MEM('o065754, 16'o000000);
`MEM('o065756, 16'o000000);
`MEM('o065760, 16'o000000);
`MEM('o065762, 16'o000000);
`MEM('o065764, 16'o000000);
`MEM('o065766, 16'o000000);
`MEM('o065770, 16'o000000);
`MEM('o065772, 16'o000000);
`MEM('o065774, 16'o000000);
`MEM('o065776, 16'o000000);
`MEM('o066000, 16'o000000);
`MEM('o066002, 16'o000000);
`MEM('o066004, 16'o000000);
`MEM('o066006, 16'o000000);
`MEM('o066010, 16'o000000);
`MEM('o066012, 16'o000000);
`MEM('o066014, 16'o000000);
`MEM('o066016, 16'o000000);
`MEM('o066020, 16'o000000);
`MEM('o066022, 16'o000000);
`MEM('o066024, 16'o000000);
`MEM('o066026, 16'o000000);
`MEM('o066030, 16'o000000);
`MEM('o066032, 16'o000000);
`MEM('o066034, 16'o000000);
`MEM('o066036, 16'o000000);
`MEM('o066040, 16'o000000);
`MEM('o066042, 16'o000000);
`MEM('o066044, 16'o000000);
`MEM('o066046, 16'o000000);
`MEM('o066050, 16'o000000);
`MEM('o066052, 16'o000000);
`MEM('o066054, 16'o000000);
`MEM('o066056, 16'o000000);
`MEM('o066060, 16'o000000);
`MEM('o066062, 16'o000000);
`MEM('o066064, 16'o000000);
`MEM('o066066, 16'o000000);
`MEM('o066070, 16'o000000);
`MEM('o066072, 16'o000000);
`MEM('o066074, 16'o000000);
`MEM('o066076, 16'o000000);
`MEM('o066100, 16'o000000);
`MEM('o066102, 16'o000000);
`MEM('o066104, 16'o000000);
`MEM('o066106, 16'o000000);
`MEM('o066110, 16'o000000);
`MEM('o066112, 16'o000000);
`MEM('o066114, 16'o000000);
`MEM('o066116, 16'o000000);
`MEM('o066120, 16'o000000);
`MEM('o066122, 16'o000000);
`MEM('o066124, 16'o000000);
`MEM('o066126, 16'o000000);
`MEM('o066130, 16'o000000);
`MEM('o066132, 16'o000000);
`MEM('o066134, 16'o000000);
`MEM('o066136, 16'o000000);
`MEM('o066140, 16'o000000);
`MEM('o066142, 16'o000000);
`MEM('o066144, 16'o000000);
`MEM('o066146, 16'o000000);
`MEM('o066150, 16'o000000);
`MEM('o066152, 16'o000000);
`MEM('o066154, 16'o000000);
`MEM('o066156, 16'o000000);
`MEM('o066160, 16'o000000);
`MEM('o066162, 16'o000000);
`MEM('o066164, 16'o000000);
`MEM('o066166, 16'o000000);
`MEM('o066170, 16'o000000);
`MEM('o066172, 16'o000000);
`MEM('o066174, 16'o000000);
`MEM('o066176, 16'o000000);
`MEM('o066200, 16'o000000);
`MEM('o066202, 16'o000000);
`MEM('o066204, 16'o000000);
`MEM('o066206, 16'o000000);
`MEM('o066210, 16'o000000);
`MEM('o066212, 16'o000000);
`MEM('o066214, 16'o000000);
`MEM('o066216, 16'o000000);
`MEM('o066220, 16'o000000);
`MEM('o066222, 16'o000000);
`MEM('o066224, 16'o000000);
`MEM('o066226, 16'o000000);
`MEM('o066230, 16'o000000);
`MEM('o066232, 16'o000000);
`MEM('o066234, 16'o000000);
`MEM('o066236, 16'o000000);
`MEM('o066240, 16'o000000);
`MEM('o066242, 16'o000000);
`MEM('o066244, 16'o000000);
`MEM('o066246, 16'o000000);
`MEM('o066250, 16'o000000);
`MEM('o066252, 16'o000000);
`MEM('o066254, 16'o000000);
`MEM('o066256, 16'o000000);
`MEM('o066260, 16'o000000);
`MEM('o066262, 16'o000000);
`MEM('o066264, 16'o000000);
`MEM('o066266, 16'o000000);
`MEM('o066270, 16'o000000);
`MEM('o066272, 16'o000000);
`MEM('o066274, 16'o000000);
`MEM('o066276, 16'o000000);
`MEM('o066300, 16'o000000);
`MEM('o066302, 16'o000000);
`MEM('o066304, 16'o000000);
`MEM('o066306, 16'o000000);
`MEM('o066310, 16'o000000);
`MEM('o066312, 16'o000000);
`MEM('o066314, 16'o000000);
`MEM('o066316, 16'o000000);
`MEM('o066320, 16'o000000);
`MEM('o066322, 16'o000000);
`MEM('o066324, 16'o000000);
`MEM('o066326, 16'o000000);
`MEM('o066330, 16'o000000);
`MEM('o066332, 16'o000000);
`MEM('o066334, 16'o000000);
`MEM('o066336, 16'o000000);
`MEM('o066340, 16'o000000);
`MEM('o066342, 16'o000000);
`MEM('o066344, 16'o000000);
`MEM('o066346, 16'o000000);
`MEM('o066350, 16'o000000);
`MEM('o066352, 16'o000000);
`MEM('o066354, 16'o000000);
`MEM('o066356, 16'o000000);
`MEM('o066360, 16'o000000);
`MEM('o066362, 16'o000000);
`MEM('o066364, 16'o000000);
`MEM('o066366, 16'o000000);
`MEM('o066370, 16'o000000);
`MEM('o066372, 16'o000000);
`MEM('o066374, 16'o000000);
`MEM('o066376, 16'o000000);
`MEM('o066400, 16'o000000);
`MEM('o066402, 16'o000000);
`MEM('o066404, 16'o000000);
`MEM('o066406, 16'o000000);
`MEM('o066410, 16'o000000);
`MEM('o066412, 16'o000000);
`MEM('o066414, 16'o000000);
`MEM('o066416, 16'o000000);
`MEM('o066420, 16'o000000);
`MEM('o066422, 16'o000000);
`MEM('o066424, 16'o000000);
`MEM('o066426, 16'o000000);
`MEM('o066430, 16'o000000);
`MEM('o066432, 16'o000000);
`MEM('o066434, 16'o000000);
`MEM('o066436, 16'o000000);
`MEM('o066440, 16'o000000);
`MEM('o066442, 16'o000000);
`MEM('o066444, 16'o000000);
`MEM('o066446, 16'o000000);
`MEM('o066450, 16'o000000);
`MEM('o066452, 16'o000000);
`MEM('o066454, 16'o000000);
`MEM('o066456, 16'o000000);
`MEM('o066460, 16'o000000);
`MEM('o066462, 16'o000000);
`MEM('o066464, 16'o000000);
`MEM('o066466, 16'o000000);
`MEM('o066470, 16'o000000);
`MEM('o066472, 16'o000000);
`MEM('o066474, 16'o000000);
`MEM('o066476, 16'o000000);
`MEM('o066500, 16'o000000);
`MEM('o066502, 16'o000000);
`MEM('o066504, 16'o000000);
`MEM('o066506, 16'o000000);
`MEM('o066510, 16'o000000);
`MEM('o066512, 16'o000000);
`MEM('o066514, 16'o000000);
`MEM('o066516, 16'o000000);
`MEM('o066520, 16'o000000);
`MEM('o066522, 16'o000000);
`MEM('o066524, 16'o000000);
`MEM('o066526, 16'o000000);
`MEM('o066530, 16'o000000);
`MEM('o066532, 16'o000000);
`MEM('o066534, 16'o000000);
`MEM('o066536, 16'o000000);
`MEM('o066540, 16'o000000);
`MEM('o066542, 16'o000000);
`MEM('o066544, 16'o000000);
`MEM('o066546, 16'o000000);
`MEM('o066550, 16'o000000);
`MEM('o066552, 16'o000000);
`MEM('o066554, 16'o000000);
`MEM('o066556, 16'o000000);
`MEM('o066560, 16'o000000);
`MEM('o066562, 16'o000000);
`MEM('o066564, 16'o000000);
`MEM('o066566, 16'o000000);
`MEM('o066570, 16'o000000);
`MEM('o066572, 16'o000000);
`MEM('o066574, 16'o000000);
`MEM('o066576, 16'o000000);
`MEM('o066600, 16'o000000);
`MEM('o066602, 16'o000000);
`MEM('o066604, 16'o000000);
`MEM('o066606, 16'o000000);
`MEM('o066610, 16'o000000);
`MEM('o066612, 16'o000000);
`MEM('o066614, 16'o000000);
`MEM('o066616, 16'o000000);
`MEM('o066620, 16'o000000);
`MEM('o066622, 16'o000000);
`MEM('o066624, 16'o000000);
`MEM('o066626, 16'o000000);
`MEM('o066630, 16'o000000);
`MEM('o066632, 16'o000000);
`MEM('o066634, 16'o000000);
`MEM('o066636, 16'o000000);
`MEM('o066640, 16'o000000);
`MEM('o066642, 16'o000000);
`MEM('o066644, 16'o000000);
`MEM('o066646, 16'o000000);
`MEM('o066650, 16'o000000);
`MEM('o066652, 16'o000000);
`MEM('o066654, 16'o000000);
`MEM('o066656, 16'o000000);
`MEM('o066660, 16'o000000);
`MEM('o066662, 16'o000000);
`MEM('o066664, 16'o000000);
`MEM('o066666, 16'o000000);
`MEM('o066670, 16'o000000);
`MEM('o066672, 16'o000000);
`MEM('o066674, 16'o000000);
`MEM('o066676, 16'o000000);
`MEM('o066700, 16'o000000);
`MEM('o066702, 16'o000000);
`MEM('o066704, 16'o000000);
`MEM('o066706, 16'o000000);
`MEM('o066710, 16'o000000);
`MEM('o066712, 16'o000000);
`MEM('o066714, 16'o000000);
`MEM('o066716, 16'o000000);
`MEM('o066720, 16'o000000);
`MEM('o066722, 16'o000000);
`MEM('o066724, 16'o000000);
`MEM('o066726, 16'o000000);
`MEM('o066730, 16'o000000);
`MEM('o066732, 16'o000000);
`MEM('o066734, 16'o000000);
`MEM('o066736, 16'o000000);
`MEM('o066740, 16'o000000);
`MEM('o066742, 16'o000000);
`MEM('o066744, 16'o000000);
`MEM('o066746, 16'o000000);
`MEM('o066750, 16'o000000);
`MEM('o066752, 16'o000000);
`MEM('o066754, 16'o000000);
`MEM('o066756, 16'o000000);
`MEM('o066760, 16'o000000);
`MEM('o066762, 16'o000000);
`MEM('o066764, 16'o000000);
`MEM('o066766, 16'o000000);
`MEM('o066770, 16'o000000);
`MEM('o066772, 16'o000000);
`MEM('o066774, 16'o000000);
`MEM('o066776, 16'o000000);
`MEM('o067000, 16'o000000);
`MEM('o067002, 16'o000000);
`MEM('o067004, 16'o000000);
`MEM('o067006, 16'o000000);
`MEM('o067010, 16'o000000);
`MEM('o067012, 16'o000000);
`MEM('o067014, 16'o000000);
`MEM('o067016, 16'o000000);
`MEM('o067020, 16'o000000);
`MEM('o067022, 16'o000000);
`MEM('o067024, 16'o000000);
`MEM('o067026, 16'o000000);
`MEM('o067030, 16'o000000);
`MEM('o067032, 16'o000000);
`MEM('o067034, 16'o000000);
`MEM('o067036, 16'o000000);
`MEM('o067040, 16'o000000);
`MEM('o067042, 16'o000000);
`MEM('o067044, 16'o000000);
`MEM('o067046, 16'o000000);
`MEM('o067050, 16'o000000);
`MEM('o067052, 16'o000000);
`MEM('o067054, 16'o000000);
`MEM('o067056, 16'o000000);
`MEM('o067060, 16'o000000);
`MEM('o067062, 16'o000000);
`MEM('o067064, 16'o000000);
`MEM('o067066, 16'o000000);
`MEM('o067070, 16'o000000);
`MEM('o067072, 16'o000000);
`MEM('o067074, 16'o000000);
`MEM('o067076, 16'o000000);
`MEM('o067100, 16'o000000);
`MEM('o067102, 16'o000000);
`MEM('o067104, 16'o000000);
`MEM('o067106, 16'o000000);
`MEM('o067110, 16'o000000);
`MEM('o067112, 16'o000000);
`MEM('o067114, 16'o000000);
`MEM('o067116, 16'o000000);
`MEM('o067120, 16'o000000);
`MEM('o067122, 16'o000000);
`MEM('o067124, 16'o000000);
`MEM('o067126, 16'o000000);
`MEM('o067130, 16'o000000);
`MEM('o067132, 16'o000000);
`MEM('o067134, 16'o000000);
`MEM('o067136, 16'o000000);
`MEM('o067140, 16'o000000);
`MEM('o067142, 16'o000000);
`MEM('o067144, 16'o000000);
`MEM('o067146, 16'o000000);
`MEM('o067150, 16'o000000);
`MEM('o067152, 16'o000000);
`MEM('o067154, 16'o000000);
`MEM('o067156, 16'o000000);
`MEM('o067160, 16'o000000);
`MEM('o067162, 16'o000000);
`MEM('o067164, 16'o000000);
`MEM('o067166, 16'o000000);
`MEM('o067170, 16'o000000);
`MEM('o067172, 16'o000000);
`MEM('o067174, 16'o000000);
`MEM('o067176, 16'o000000);
`MEM('o067200, 16'o000000);
`MEM('o067202, 16'o000000);
`MEM('o067204, 16'o000000);
`MEM('o067206, 16'o000000);
`MEM('o067210, 16'o000000);
`MEM('o067212, 16'o000000);
`MEM('o067214, 16'o000000);
`MEM('o067216, 16'o000000);
`MEM('o067220, 16'o000000);
`MEM('o067222, 16'o000000);
`MEM('o067224, 16'o000000);
`MEM('o067226, 16'o000000);
`MEM('o067230, 16'o000000);
`MEM('o067232, 16'o000000);
`MEM('o067234, 16'o000000);
`MEM('o067236, 16'o000000);
`MEM('o067240, 16'o000000);
`MEM('o067242, 16'o000000);
`MEM('o067244, 16'o000000);
`MEM('o067246, 16'o000000);
`MEM('o067250, 16'o000000);
`MEM('o067252, 16'o000000);
`MEM('o067254, 16'o000000);
`MEM('o067256, 16'o000000);
`MEM('o067260, 16'o000000);
`MEM('o067262, 16'o000000);
`MEM('o067264, 16'o000000);
`MEM('o067266, 16'o000000);
`MEM('o067270, 16'o000000);
`MEM('o067272, 16'o000000);
`MEM('o067274, 16'o000000);
`MEM('o067276, 16'o000000);
`MEM('o067300, 16'o000000);
`MEM('o067302, 16'o000000);
`MEM('o067304, 16'o000000);
`MEM('o067306, 16'o000000);
`MEM('o067310, 16'o000000);
`MEM('o067312, 16'o000000);
`MEM('o067314, 16'o000000);
`MEM('o067316, 16'o000000);
`MEM('o067320, 16'o000000);
`MEM('o067322, 16'o000000);
`MEM('o067324, 16'o000000);
`MEM('o067326, 16'o000000);
`MEM('o067330, 16'o000000);
`MEM('o067332, 16'o000000);
`MEM('o067334, 16'o000000);
`MEM('o067336, 16'o000000);
`MEM('o067340, 16'o000000);
`MEM('o067342, 16'o000000);
`MEM('o067344, 16'o000000);
`MEM('o067346, 16'o000000);
`MEM('o067350, 16'o000000);
`MEM('o067352, 16'o000000);
`MEM('o067354, 16'o000000);
`MEM('o067356, 16'o000000);
`MEM('o067360, 16'o000000);
`MEM('o067362, 16'o000000);
`MEM('o067364, 16'o000000);
`MEM('o067366, 16'o000000);
`MEM('o067370, 16'o000000);
`MEM('o067372, 16'o000000);
`MEM('o067374, 16'o000000);
`MEM('o067376, 16'o000000);
`MEM('o067400, 16'o000000);
`MEM('o067402, 16'o000000);
`MEM('o067404, 16'o000000);
`MEM('o067406, 16'o000000);
`MEM('o067410, 16'o000000);
`MEM('o067412, 16'o000000);
`MEM('o067414, 16'o000000);
`MEM('o067416, 16'o000000);
`MEM('o067420, 16'o000000);
`MEM('o067422, 16'o000000);
`MEM('o067424, 16'o000000);
`MEM('o067426, 16'o000000);
`MEM('o067430, 16'o000000);
`MEM('o067432, 16'o000000);
`MEM('o067434, 16'o000000);
`MEM('o067436, 16'o000000);
`MEM('o067440, 16'o000000);
`MEM('o067442, 16'o000000);
`MEM('o067444, 16'o000000);
`MEM('o067446, 16'o000000);
`MEM('o067450, 16'o000000);
`MEM('o067452, 16'o000000);
`MEM('o067454, 16'o000000);
`MEM('o067456, 16'o000000);
`MEM('o067460, 16'o000000);
`MEM('o067462, 16'o000000);
`MEM('o067464, 16'o000000);
`MEM('o067466, 16'o000000);
`MEM('o067470, 16'o000000);
`MEM('o067472, 16'o000000);
`MEM('o067474, 16'o000000);
`MEM('o067476, 16'o000000);
`MEM('o067500, 16'o000000);
`MEM('o067502, 16'o000000);
`MEM('o067504, 16'o000000);
`MEM('o067506, 16'o000000);
`MEM('o067510, 16'o000000);
`MEM('o067512, 16'o000000);
`MEM('o067514, 16'o000000);
`MEM('o067516, 16'o000000);
`MEM('o067520, 16'o000000);
`MEM('o067522, 16'o000000);
`MEM('o067524, 16'o000000);
`MEM('o067526, 16'o000000);
`MEM('o067530, 16'o000000);
`MEM('o067532, 16'o000000);
`MEM('o067534, 16'o000000);
`MEM('o067536, 16'o000000);
`MEM('o067540, 16'o000000);
`MEM('o067542, 16'o000000);
`MEM('o067544, 16'o000000);
`MEM('o067546, 16'o000000);
`MEM('o067550, 16'o000000);
`MEM('o067552, 16'o000000);
`MEM('o067554, 16'o000000);
`MEM('o067556, 16'o000000);
`MEM('o067560, 16'o000000);
`MEM('o067562, 16'o000000);
`MEM('o067564, 16'o000000);
`MEM('o067566, 16'o000000);
`MEM('o067570, 16'o000000);
`MEM('o067572, 16'o000000);
`MEM('o067574, 16'o000000);
`MEM('o067576, 16'o000000);
`MEM('o067600, 16'o000000);
`MEM('o067602, 16'o000000);
`MEM('o067604, 16'o000000);
`MEM('o067606, 16'o000000);
`MEM('o067610, 16'o000000);
`MEM('o067612, 16'o000000);
`MEM('o067614, 16'o000000);
`MEM('o067616, 16'o000000);
`MEM('o067620, 16'o000000);
`MEM('o067622, 16'o000000);
`MEM('o067624, 16'o000000);
`MEM('o067626, 16'o000000);
`MEM('o067630, 16'o000000);
`MEM('o067632, 16'o000000);
`MEM('o067634, 16'o000000);
`MEM('o067636, 16'o000000);
`MEM('o067640, 16'o000000);
`MEM('o067642, 16'o000000);
`MEM('o067644, 16'o000000);
`MEM('o067646, 16'o000000);
`MEM('o067650, 16'o000000);
`MEM('o067652, 16'o000000);
`MEM('o067654, 16'o000000);
`MEM('o067656, 16'o000000);
`MEM('o067660, 16'o000000);
`MEM('o067662, 16'o000000);
`MEM('o067664, 16'o000000);
`MEM('o067666, 16'o000000);
`MEM('o067670, 16'o000000);
`MEM('o067672, 16'o000000);
`MEM('o067674, 16'o000000);
`MEM('o067676, 16'o000000);
`MEM('o067700, 16'o000000);
`MEM('o067702, 16'o000000);
`MEM('o067704, 16'o000000);
`MEM('o067706, 16'o000000);
`MEM('o067710, 16'o000000);
`MEM('o067712, 16'o000000);
`MEM('o067714, 16'o000000);
`MEM('o067716, 16'o000000);
`MEM('o067720, 16'o000000);
`MEM('o067722, 16'o000000);
`MEM('o067724, 16'o000000);
`MEM('o067726, 16'o000000);
`MEM('o067730, 16'o000000);
`MEM('o067732, 16'o000000);
`MEM('o067734, 16'o000000);
`MEM('o067736, 16'o000000);
`MEM('o067740, 16'o000000);
`MEM('o067742, 16'o000000);
`MEM('o067744, 16'o000000);
`MEM('o067746, 16'o000000);
`MEM('o067750, 16'o000000);
`MEM('o067752, 16'o000000);
`MEM('o067754, 16'o000000);
`MEM('o067756, 16'o000000);
`MEM('o067760, 16'o000000);
`MEM('o067762, 16'o000000);
`MEM('o067764, 16'o000000);
`MEM('o067766, 16'o000000);
`MEM('o067770, 16'o000000);
`MEM('o067772, 16'o000000);
`MEM('o067774, 16'o000000);
`MEM('o067776, 16'o000000);
`MEM('o070000, 16'o000000);
`MEM('o070002, 16'o000000);
`MEM('o070004, 16'o000000);
`MEM('o070006, 16'o000000);
`MEM('o070010, 16'o000000);
`MEM('o070012, 16'o000000);
`MEM('o070014, 16'o000000);
`MEM('o070016, 16'o000000);
`MEM('o070020, 16'o000000);
`MEM('o070022, 16'o000000);
`MEM('o070024, 16'o000000);
`MEM('o070026, 16'o000000);
`MEM('o070030, 16'o000000);
`MEM('o070032, 16'o000000);
`MEM('o070034, 16'o000000);
`MEM('o070036, 16'o000000);
`MEM('o070040, 16'o000000);
`MEM('o070042, 16'o000000);
`MEM('o070044, 16'o000000);
`MEM('o070046, 16'o000000);
`MEM('o070050, 16'o000000);
`MEM('o070052, 16'o000000);
`MEM('o070054, 16'o000000);
`MEM('o070056, 16'o000000);
`MEM('o070060, 16'o000000);
`MEM('o070062, 16'o000000);
`MEM('o070064, 16'o000000);
`MEM('o070066, 16'o000000);
`MEM('o070070, 16'o000000);
`MEM('o070072, 16'o000000);
`MEM('o070074, 16'o000000);
`MEM('o070076, 16'o000000);
`MEM('o070100, 16'o000000);
`MEM('o070102, 16'o000000);
`MEM('o070104, 16'o000000);
`MEM('o070106, 16'o000000);
`MEM('o070110, 16'o000000);
`MEM('o070112, 16'o000000);
`MEM('o070114, 16'o000000);
`MEM('o070116, 16'o000000);
`MEM('o070120, 16'o000000);
`MEM('o070122, 16'o000000);
`MEM('o070124, 16'o000000);
`MEM('o070126, 16'o000000);
`MEM('o070130, 16'o000000);
`MEM('o070132, 16'o000000);
`MEM('o070134, 16'o000000);
`MEM('o070136, 16'o000000);
`MEM('o070140, 16'o000000);
`MEM('o070142, 16'o000000);
`MEM('o070144, 16'o000000);
`MEM('o070146, 16'o000000);
`MEM('o070150, 16'o000000);
`MEM('o070152, 16'o000000);
`MEM('o070154, 16'o000000);
`MEM('o070156, 16'o000000);
`MEM('o070160, 16'o000000);
`MEM('o070162, 16'o000000);
`MEM('o070164, 16'o000000);
`MEM('o070166, 16'o000000);
`MEM('o070170, 16'o000000);
`MEM('o070172, 16'o000000);
`MEM('o070174, 16'o000000);
`MEM('o070176, 16'o000000);
`MEM('o070200, 16'o000000);
`MEM('o070202, 16'o000000);
`MEM('o070204, 16'o000000);
`MEM('o070206, 16'o000000);
`MEM('o070210, 16'o000000);
`MEM('o070212, 16'o000000);
`MEM('o070214, 16'o000000);
`MEM('o070216, 16'o000000);
`MEM('o070220, 16'o000000);
`MEM('o070222, 16'o000000);
`MEM('o070224, 16'o000000);
`MEM('o070226, 16'o000000);
`MEM('o070230, 16'o000000);
`MEM('o070232, 16'o000000);
`MEM('o070234, 16'o000000);
`MEM('o070236, 16'o000000);
`MEM('o070240, 16'o000000);
`MEM('o070242, 16'o000000);
`MEM('o070244, 16'o000000);
`MEM('o070246, 16'o000000);
`MEM('o070250, 16'o000000);
`MEM('o070252, 16'o000000);
`MEM('o070254, 16'o000000);
`MEM('o070256, 16'o000000);
`MEM('o070260, 16'o000000);
`MEM('o070262, 16'o000000);
`MEM('o070264, 16'o000000);
`MEM('o070266, 16'o000000);
`MEM('o070270, 16'o000000);
`MEM('o070272, 16'o000000);
`MEM('o070274, 16'o000000);
`MEM('o070276, 16'o000000);
`MEM('o070300, 16'o000000);
`MEM('o070302, 16'o000000);
`MEM('o070304, 16'o000000);
`MEM('o070306, 16'o000000);
`MEM('o070310, 16'o000000);
`MEM('o070312, 16'o000000);
`MEM('o070314, 16'o000000);
`MEM('o070316, 16'o000000);
`MEM('o070320, 16'o000000);
`MEM('o070322, 16'o000000);
`MEM('o070324, 16'o000000);
`MEM('o070326, 16'o000000);
`MEM('o070330, 16'o000000);
`MEM('o070332, 16'o000000);
`MEM('o070334, 16'o000000);
`MEM('o070336, 16'o000000);
`MEM('o070340, 16'o000000);
`MEM('o070342, 16'o000000);
`MEM('o070344, 16'o000000);
`MEM('o070346, 16'o000000);
`MEM('o070350, 16'o000000);
`MEM('o070352, 16'o000000);
`MEM('o070354, 16'o000000);
`MEM('o070356, 16'o000000);
`MEM('o070360, 16'o000000);
`MEM('o070362, 16'o000000);
`MEM('o070364, 16'o000000);
`MEM('o070366, 16'o000000);
`MEM('o070370, 16'o000000);
`MEM('o070372, 16'o000000);
`MEM('o070374, 16'o000000);
`MEM('o070376, 16'o000000);
`MEM('o070400, 16'o000000);
`MEM('o070402, 16'o000000);
`MEM('o070404, 16'o000000);
`MEM('o070406, 16'o000000);
`MEM('o070410, 16'o000000);
`MEM('o070412, 16'o000000);
`MEM('o070414, 16'o000000);
`MEM('o070416, 16'o000000);
`MEM('o070420, 16'o000000);
`MEM('o070422, 16'o000000);
`MEM('o070424, 16'o000000);
`MEM('o070426, 16'o000000);
`MEM('o070430, 16'o000000);
`MEM('o070432, 16'o000000);
`MEM('o070434, 16'o000000);
`MEM('o070436, 16'o000000);
`MEM('o070440, 16'o000000);
`MEM('o070442, 16'o000000);
`MEM('o070444, 16'o000000);
`MEM('o070446, 16'o000000);
`MEM('o070450, 16'o000000);
`MEM('o070452, 16'o000000);
`MEM('o070454, 16'o000000);
`MEM('o070456, 16'o000000);
`MEM('o070460, 16'o000000);
`MEM('o070462, 16'o000000);
`MEM('o070464, 16'o000000);
`MEM('o070466, 16'o000000);
`MEM('o070470, 16'o000000);
`MEM('o070472, 16'o000000);
`MEM('o070474, 16'o000000);
`MEM('o070476, 16'o000000);
`MEM('o070500, 16'o000000);
`MEM('o070502, 16'o000000);
`MEM('o070504, 16'o000000);
`MEM('o070506, 16'o000000);
`MEM('o070510, 16'o000000);
`MEM('o070512, 16'o000000);
`MEM('o070514, 16'o000000);
`MEM('o070516, 16'o000000);
`MEM('o070520, 16'o000000);
`MEM('o070522, 16'o000000);
`MEM('o070524, 16'o000000);
`MEM('o070526, 16'o000000);
`MEM('o070530, 16'o000000);
`MEM('o070532, 16'o000000);
`MEM('o070534, 16'o000000);
`MEM('o070536, 16'o000000);
`MEM('o070540, 16'o000000);
`MEM('o070542, 16'o000000);
`MEM('o070544, 16'o000000);
`MEM('o070546, 16'o000000);
`MEM('o070550, 16'o000000);
`MEM('o070552, 16'o000000);
`MEM('o070554, 16'o000000);
`MEM('o070556, 16'o000000);
`MEM('o070560, 16'o000000);
`MEM('o070562, 16'o000000);
`MEM('o070564, 16'o000000);
`MEM('o070566, 16'o000000);
`MEM('o070570, 16'o000000);
`MEM('o070572, 16'o000000);
`MEM('o070574, 16'o000000);
`MEM('o070576, 16'o000000);
`MEM('o070600, 16'o000000);
`MEM('o070602, 16'o000000);
`MEM('o070604, 16'o000000);
`MEM('o070606, 16'o000000);
`MEM('o070610, 16'o000000);
`MEM('o070612, 16'o000000);
`MEM('o070614, 16'o000000);
`MEM('o070616, 16'o000000);
`MEM('o070620, 16'o000000);
`MEM('o070622, 16'o000000);
`MEM('o070624, 16'o000000);
`MEM('o070626, 16'o000000);
`MEM('o070630, 16'o000000);
`MEM('o070632, 16'o000000);
`MEM('o070634, 16'o000000);
`MEM('o070636, 16'o000000);
`MEM('o070640, 16'o000000);
`MEM('o070642, 16'o000000);
`MEM('o070644, 16'o000000);
`MEM('o070646, 16'o000000);
`MEM('o070650, 16'o000000);
`MEM('o070652, 16'o000000);
`MEM('o070654, 16'o000000);
`MEM('o070656, 16'o000000);
`MEM('o070660, 16'o000000);
`MEM('o070662, 16'o000000);
`MEM('o070664, 16'o000000);
`MEM('o070666, 16'o000000);
`MEM('o070670, 16'o000000);
`MEM('o070672, 16'o000000);
`MEM('o070674, 16'o000000);
`MEM('o070676, 16'o000000);
`MEM('o070700, 16'o000000);
`MEM('o070702, 16'o000000);
`MEM('o070704, 16'o000000);
`MEM('o070706, 16'o000000);
`MEM('o070710, 16'o000000);
`MEM('o070712, 16'o000000);
`MEM('o070714, 16'o000000);
`MEM('o070716, 16'o000000);
`MEM('o070720, 16'o000000);
`MEM('o070722, 16'o000000);
`MEM('o070724, 16'o000000);
`MEM('o070726, 16'o000000);
`MEM('o070730, 16'o000000);
`MEM('o070732, 16'o000000);
`MEM('o070734, 16'o000000);
`MEM('o070736, 16'o000000);
`MEM('o070740, 16'o000000);
`MEM('o070742, 16'o000000);
`MEM('o070744, 16'o000000);
`MEM('o070746, 16'o000000);
`MEM('o070750, 16'o000000);
`MEM('o070752, 16'o000000);
`MEM('o070754, 16'o000000);
`MEM('o070756, 16'o000000);
`MEM('o070760, 16'o000000);
`MEM('o070762, 16'o000000);
`MEM('o070764, 16'o000000);
`MEM('o070766, 16'o000000);
`MEM('o070770, 16'o000000);
`MEM('o070772, 16'o000000);
`MEM('o070774, 16'o000000);
`MEM('o070776, 16'o000000);
`MEM('o071000, 16'o000000);
`MEM('o071002, 16'o000000);
`MEM('o071004, 16'o000000);
`MEM('o071006, 16'o000000);
`MEM('o071010, 16'o000000);
`MEM('o071012, 16'o000000);
`MEM('o071014, 16'o000000);
`MEM('o071016, 16'o000000);
`MEM('o071020, 16'o000000);
`MEM('o071022, 16'o000000);
`MEM('o071024, 16'o000000);
`MEM('o071026, 16'o000000);
`MEM('o071030, 16'o000000);
`MEM('o071032, 16'o000000);
`MEM('o071034, 16'o000000);
`MEM('o071036, 16'o000000);
`MEM('o071040, 16'o000000);
`MEM('o071042, 16'o000000);
`MEM('o071044, 16'o000000);
`MEM('o071046, 16'o000000);
`MEM('o071050, 16'o000000);
`MEM('o071052, 16'o000000);
`MEM('o071054, 16'o000000);
`MEM('o071056, 16'o000000);
`MEM('o071060, 16'o000000);
`MEM('o071062, 16'o000000);
`MEM('o071064, 16'o000000);
`MEM('o071066, 16'o000000);
`MEM('o071070, 16'o000000);
`MEM('o071072, 16'o000000);
`MEM('o071074, 16'o000000);
`MEM('o071076, 16'o000000);
`MEM('o071100, 16'o000000);
`MEM('o071102, 16'o000000);
`MEM('o071104, 16'o000000);
`MEM('o071106, 16'o000000);
`MEM('o071110, 16'o000000);
`MEM('o071112, 16'o000000);
`MEM('o071114, 16'o000000);
`MEM('o071116, 16'o000000);
`MEM('o071120, 16'o000000);
`MEM('o071122, 16'o000000);
`MEM('o071124, 16'o000000);
`MEM('o071126, 16'o000000);
`MEM('o071130, 16'o000000);
`MEM('o071132, 16'o000000);
`MEM('o071134, 16'o000000);
`MEM('o071136, 16'o000000);
`MEM('o071140, 16'o000000);
`MEM('o071142, 16'o000000);
`MEM('o071144, 16'o000000);
`MEM('o071146, 16'o000000);
`MEM('o071150, 16'o000000);
`MEM('o071152, 16'o000000);
`MEM('o071154, 16'o000000);
`MEM('o071156, 16'o000000);
`MEM('o071160, 16'o000000);
`MEM('o071162, 16'o000000);
`MEM('o071164, 16'o000000);
`MEM('o071166, 16'o000000);
`MEM('o071170, 16'o000000);
`MEM('o071172, 16'o000000);
`MEM('o071174, 16'o000000);
`MEM('o071176, 16'o000000);
`MEM('o071200, 16'o000000);
`MEM('o071202, 16'o000000);
`MEM('o071204, 16'o000000);
`MEM('o071206, 16'o000000);
`MEM('o071210, 16'o000000);
`MEM('o071212, 16'o000000);
`MEM('o071214, 16'o000000);
`MEM('o071216, 16'o000000);
`MEM('o071220, 16'o000000);
`MEM('o071222, 16'o000000);
`MEM('o071224, 16'o000000);
`MEM('o071226, 16'o000000);
`MEM('o071230, 16'o000000);
`MEM('o071232, 16'o000000);
`MEM('o071234, 16'o000000);
`MEM('o071236, 16'o000000);
`MEM('o071240, 16'o000000);
`MEM('o071242, 16'o000000);
`MEM('o071244, 16'o000000);
`MEM('o071246, 16'o000000);
`MEM('o071250, 16'o000000);
`MEM('o071252, 16'o000000);
`MEM('o071254, 16'o000000);
`MEM('o071256, 16'o000000);
`MEM('o071260, 16'o000000);
`MEM('o071262, 16'o000000);
`MEM('o071264, 16'o000000);
`MEM('o071266, 16'o000000);
`MEM('o071270, 16'o000000);
`MEM('o071272, 16'o000000);
`MEM('o071274, 16'o000000);
`MEM('o071276, 16'o000000);
`MEM('o071300, 16'o000000);
`MEM('o071302, 16'o000000);
`MEM('o071304, 16'o000000);
`MEM('o071306, 16'o000000);
`MEM('o071310, 16'o000000);
`MEM('o071312, 16'o000000);
`MEM('o071314, 16'o000000);
`MEM('o071316, 16'o000000);
`MEM('o071320, 16'o000000);
`MEM('o071322, 16'o000000);
`MEM('o071324, 16'o000000);
`MEM('o071326, 16'o000000);
`MEM('o071330, 16'o000000);
`MEM('o071332, 16'o000000);
`MEM('o071334, 16'o000000);
`MEM('o071336, 16'o000000);
`MEM('o071340, 16'o000000);
`MEM('o071342, 16'o000000);
`MEM('o071344, 16'o000000);
`MEM('o071346, 16'o000000);
`MEM('o071350, 16'o000000);
`MEM('o071352, 16'o000000);
`MEM('o071354, 16'o000000);
`MEM('o071356, 16'o000000);
`MEM('o071360, 16'o000000);
`MEM('o071362, 16'o000000);
`MEM('o071364, 16'o000000);
`MEM('o071366, 16'o000000);
`MEM('o071370, 16'o000000);
`MEM('o071372, 16'o000000);
`MEM('o071374, 16'o000000);
`MEM('o071376, 16'o000000);
`MEM('o071400, 16'o000000);
`MEM('o071402, 16'o000000);
`MEM('o071404, 16'o000000);
`MEM('o071406, 16'o000000);
`MEM('o071410, 16'o000000);
`MEM('o071412, 16'o000000);
`MEM('o071414, 16'o000000);
`MEM('o071416, 16'o000000);
`MEM('o071420, 16'o000000);
`MEM('o071422, 16'o000000);
`MEM('o071424, 16'o000000);
`MEM('o071426, 16'o000000);
`MEM('o071430, 16'o000000);
`MEM('o071432, 16'o000000);
`MEM('o071434, 16'o000000);
`MEM('o071436, 16'o000000);
`MEM('o071440, 16'o000000);
`MEM('o071442, 16'o000000);
`MEM('o071444, 16'o000000);
`MEM('o071446, 16'o000000);
`MEM('o071450, 16'o000000);
`MEM('o071452, 16'o000000);
`MEM('o071454, 16'o000000);
`MEM('o071456, 16'o000000);
`MEM('o071460, 16'o000000);
`MEM('o071462, 16'o000000);
`MEM('o071464, 16'o000000);
`MEM('o071466, 16'o000000);
`MEM('o071470, 16'o000000);
`MEM('o071472, 16'o000000);
`MEM('o071474, 16'o000000);
`MEM('o071476, 16'o000000);
`MEM('o071500, 16'o000000);
`MEM('o071502, 16'o000000);
`MEM('o071504, 16'o000000);
`MEM('o071506, 16'o000000);
`MEM('o071510, 16'o000000);
`MEM('o071512, 16'o000000);
`MEM('o071514, 16'o000000);
`MEM('o071516, 16'o000000);
`MEM('o071520, 16'o000000);
`MEM('o071522, 16'o000000);
`MEM('o071524, 16'o000000);
`MEM('o071526, 16'o000000);
`MEM('o071530, 16'o000000);
`MEM('o071532, 16'o000000);
`MEM('o071534, 16'o000000);
`MEM('o071536, 16'o000000);
`MEM('o071540, 16'o000000);
`MEM('o071542, 16'o000000);
`MEM('o071544, 16'o000000);
`MEM('o071546, 16'o000000);
`MEM('o071550, 16'o000000);
`MEM('o071552, 16'o000000);
`MEM('o071554, 16'o000000);
`MEM('o071556, 16'o000000);
`MEM('o071560, 16'o000000);
`MEM('o071562, 16'o000000);
`MEM('o071564, 16'o000000);
`MEM('o071566, 16'o000000);
`MEM('o071570, 16'o000000);
`MEM('o071572, 16'o000000);
`MEM('o071574, 16'o000000);
`MEM('o071576, 16'o000000);
`MEM('o071600, 16'o000000);
`MEM('o071602, 16'o000000);
`MEM('o071604, 16'o000000);
`MEM('o071606, 16'o000000);
`MEM('o071610, 16'o000000);
`MEM('o071612, 16'o000000);
`MEM('o071614, 16'o000000);
`MEM('o071616, 16'o000000);
`MEM('o071620, 16'o000000);
`MEM('o071622, 16'o000000);
`MEM('o071624, 16'o000000);
`MEM('o071626, 16'o000000);
`MEM('o071630, 16'o000000);
`MEM('o071632, 16'o000000);
`MEM('o071634, 16'o000000);
`MEM('o071636, 16'o000000);
`MEM('o071640, 16'o000000);
`MEM('o071642, 16'o000000);
`MEM('o071644, 16'o000000);
`MEM('o071646, 16'o000000);
`MEM('o071650, 16'o000000);
`MEM('o071652, 16'o000000);
`MEM('o071654, 16'o000000);
`MEM('o071656, 16'o000000);
`MEM('o071660, 16'o000000);
`MEM('o071662, 16'o000000);
`MEM('o071664, 16'o000000);
`MEM('o071666, 16'o000000);
`MEM('o071670, 16'o000000);
`MEM('o071672, 16'o000000);
`MEM('o071674, 16'o000000);
`MEM('o071676, 16'o000000);
`MEM('o071700, 16'o000000);
`MEM('o071702, 16'o000000);
`MEM('o071704, 16'o000000);
`MEM('o071706, 16'o000000);
`MEM('o071710, 16'o000000);
`MEM('o071712, 16'o000000);
`MEM('o071714, 16'o000000);
`MEM('o071716, 16'o000000);
`MEM('o071720, 16'o000000);
`MEM('o071722, 16'o000000);
`MEM('o071724, 16'o000000);
`MEM('o071726, 16'o000000);
`MEM('o071730, 16'o000000);
`MEM('o071732, 16'o000000);
`MEM('o071734, 16'o000000);
`MEM('o071736, 16'o000000);
`MEM('o071740, 16'o000000);
`MEM('o071742, 16'o000000);
`MEM('o071744, 16'o000000);
`MEM('o071746, 16'o000000);
`MEM('o071750, 16'o000000);
`MEM('o071752, 16'o000000);
`MEM('o071754, 16'o000000);
`MEM('o071756, 16'o000000);
`MEM('o071760, 16'o000000);
`MEM('o071762, 16'o000000);
`MEM('o071764, 16'o000000);
`MEM('o071766, 16'o000000);
`MEM('o071770, 16'o000000);
`MEM('o071772, 16'o000000);
`MEM('o071774, 16'o000000);
`MEM('o071776, 16'o000000);
`MEM('o072000, 16'o000000);
`MEM('o072002, 16'o000000);
`MEM('o072004, 16'o000000);
`MEM('o072006, 16'o000000);
`MEM('o072010, 16'o000000);
`MEM('o072012, 16'o000000);
`MEM('o072014, 16'o000000);
`MEM('o072016, 16'o000000);
`MEM('o072020, 16'o000000);
`MEM('o072022, 16'o000000);
`MEM('o072024, 16'o000000);
`MEM('o072026, 16'o000000);
`MEM('o072030, 16'o000000);
`MEM('o072032, 16'o000000);
`MEM('o072034, 16'o000000);
`MEM('o072036, 16'o000000);
`MEM('o072040, 16'o000000);
`MEM('o072042, 16'o000000);
`MEM('o072044, 16'o000000);
`MEM('o072046, 16'o000000);
`MEM('o072050, 16'o000000);
`MEM('o072052, 16'o000000);
`MEM('o072054, 16'o000000);
`MEM('o072056, 16'o000000);
`MEM('o072060, 16'o000000);
`MEM('o072062, 16'o000000);
`MEM('o072064, 16'o000000);
`MEM('o072066, 16'o000000);
`MEM('o072070, 16'o000000);
`MEM('o072072, 16'o000000);
`MEM('o072074, 16'o000000);
`MEM('o072076, 16'o000000);
`MEM('o072100, 16'o000000);
`MEM('o072102, 16'o000000);
`MEM('o072104, 16'o000000);
`MEM('o072106, 16'o000000);
`MEM('o072110, 16'o000000);
`MEM('o072112, 16'o000000);
`MEM('o072114, 16'o000000);
`MEM('o072116, 16'o000000);
`MEM('o072120, 16'o000000);
`MEM('o072122, 16'o000000);
`MEM('o072124, 16'o000000);
`MEM('o072126, 16'o000000);
`MEM('o072130, 16'o000000);
`MEM('o072132, 16'o000000);
`MEM('o072134, 16'o000000);
`MEM('o072136, 16'o000000);
`MEM('o072140, 16'o000000);
`MEM('o072142, 16'o000000);
`MEM('o072144, 16'o000000);
`MEM('o072146, 16'o000000);
`MEM('o072150, 16'o000000);
`MEM('o072152, 16'o000000);
`MEM('o072154, 16'o000000);
`MEM('o072156, 16'o000000);
`MEM('o072160, 16'o000000);
`MEM('o072162, 16'o000000);
`MEM('o072164, 16'o000000);
`MEM('o072166, 16'o000000);
`MEM('o072170, 16'o000000);
`MEM('o072172, 16'o000000);
`MEM('o072174, 16'o000000);
`MEM('o072176, 16'o000000);
`MEM('o072200, 16'o000000);
`MEM('o072202, 16'o000000);
`MEM('o072204, 16'o000000);
`MEM('o072206, 16'o000000);
`MEM('o072210, 16'o000000);
`MEM('o072212, 16'o000000);
`MEM('o072214, 16'o000000);
`MEM('o072216, 16'o000000);
`MEM('o072220, 16'o000000);
`MEM('o072222, 16'o000000);
`MEM('o072224, 16'o000000);
`MEM('o072226, 16'o000000);
`MEM('o072230, 16'o000000);
`MEM('o072232, 16'o000000);
`MEM('o072234, 16'o000000);
`MEM('o072236, 16'o000000);
`MEM('o072240, 16'o000000);
`MEM('o072242, 16'o000000);
`MEM('o072244, 16'o000000);
`MEM('o072246, 16'o000000);
`MEM('o072250, 16'o000000);
`MEM('o072252, 16'o000000);
`MEM('o072254, 16'o000000);
`MEM('o072256, 16'o000000);
`MEM('o072260, 16'o000000);
`MEM('o072262, 16'o000000);
`MEM('o072264, 16'o000000);
`MEM('o072266, 16'o000000);
`MEM('o072270, 16'o000000);
`MEM('o072272, 16'o000000);
`MEM('o072274, 16'o000000);
`MEM('o072276, 16'o000000);
`MEM('o072300, 16'o000000);
`MEM('o072302, 16'o000000);
`MEM('o072304, 16'o000000);
`MEM('o072306, 16'o000000);
`MEM('o072310, 16'o000000);
`MEM('o072312, 16'o000000);
`MEM('o072314, 16'o000000);
`MEM('o072316, 16'o000000);
`MEM('o072320, 16'o000000);
`MEM('o072322, 16'o000000);
`MEM('o072324, 16'o000000);
`MEM('o072326, 16'o000000);
`MEM('o072330, 16'o000000);
`MEM('o072332, 16'o000000);
`MEM('o072334, 16'o000000);
`MEM('o072336, 16'o000000);
`MEM('o072340, 16'o000000);
`MEM('o072342, 16'o000000);
`MEM('o072344, 16'o000000);
`MEM('o072346, 16'o000000);
`MEM('o072350, 16'o000000);
`MEM('o072352, 16'o000000);
`MEM('o072354, 16'o000000);
`MEM('o072356, 16'o000000);
`MEM('o072360, 16'o000000);
`MEM('o072362, 16'o000000);
`MEM('o072364, 16'o000000);
`MEM('o072366, 16'o000000);
`MEM('o072370, 16'o000000);
`MEM('o072372, 16'o000000);
`MEM('o072374, 16'o000000);
`MEM('o072376, 16'o000000);
`MEM('o072400, 16'o000000);
`MEM('o072402, 16'o000000);
`MEM('o072404, 16'o000000);
`MEM('o072406, 16'o000000);
`MEM('o072410, 16'o000000);
`MEM('o072412, 16'o000000);
`MEM('o072414, 16'o000000);
`MEM('o072416, 16'o000000);
`MEM('o072420, 16'o000000);
`MEM('o072422, 16'o000000);
`MEM('o072424, 16'o000000);
`MEM('o072426, 16'o000000);
`MEM('o072430, 16'o000000);
`MEM('o072432, 16'o000000);
`MEM('o072434, 16'o000000);
`MEM('o072436, 16'o000000);
`MEM('o072440, 16'o000000);
`MEM('o072442, 16'o000000);
`MEM('o072444, 16'o000000);
`MEM('o072446, 16'o000000);
`MEM('o072450, 16'o000000);
`MEM('o072452, 16'o000000);
`MEM('o072454, 16'o000000);
`MEM('o072456, 16'o000000);
`MEM('o072460, 16'o000000);
`MEM('o072462, 16'o000000);
`MEM('o072464, 16'o000000);
`MEM('o072466, 16'o000000);
`MEM('o072470, 16'o000000);
`MEM('o072472, 16'o000000);
`MEM('o072474, 16'o000000);
`MEM('o072476, 16'o000000);
`MEM('o072500, 16'o000000);
`MEM('o072502, 16'o000000);
`MEM('o072504, 16'o000000);
`MEM('o072506, 16'o000000);
`MEM('o072510, 16'o000000);
`MEM('o072512, 16'o000000);
`MEM('o072514, 16'o000000);
`MEM('o072516, 16'o000000);
`MEM('o072520, 16'o000000);
`MEM('o072522, 16'o000000);
`MEM('o072524, 16'o000000);
`MEM('o072526, 16'o000000);
`MEM('o072530, 16'o000000);
`MEM('o072532, 16'o000000);
`MEM('o072534, 16'o000000);
`MEM('o072536, 16'o000000);
`MEM('o072540, 16'o000000);
`MEM('o072542, 16'o000000);
`MEM('o072544, 16'o000000);
`MEM('o072546, 16'o000000);
`MEM('o072550, 16'o000000);
`MEM('o072552, 16'o000000);
`MEM('o072554, 16'o000000);
`MEM('o072556, 16'o000000);
`MEM('o072560, 16'o000000);
`MEM('o072562, 16'o000000);
`MEM('o072564, 16'o000000);
`MEM('o072566, 16'o000000);
`MEM('o072570, 16'o000000);
`MEM('o072572, 16'o000000);
`MEM('o072574, 16'o000000);
`MEM('o072576, 16'o000000);
`MEM('o072600, 16'o000000);
`MEM('o072602, 16'o000000);
`MEM('o072604, 16'o000000);
`MEM('o072606, 16'o000000);
`MEM('o072610, 16'o000000);
`MEM('o072612, 16'o000000);
`MEM('o072614, 16'o000000);
`MEM('o072616, 16'o000000);
`MEM('o072620, 16'o000000);
`MEM('o072622, 16'o000000);
`MEM('o072624, 16'o000000);
`MEM('o072626, 16'o000000);
`MEM('o072630, 16'o000000);
`MEM('o072632, 16'o000000);
`MEM('o072634, 16'o000000);
`MEM('o072636, 16'o000000);
`MEM('o072640, 16'o000000);
`MEM('o072642, 16'o000000);
`MEM('o072644, 16'o000000);
`MEM('o072646, 16'o000000);
`MEM('o072650, 16'o000000);
`MEM('o072652, 16'o000000);
`MEM('o072654, 16'o000000);
`MEM('o072656, 16'o000000);
`MEM('o072660, 16'o000000);
`MEM('o072662, 16'o000000);
`MEM('o072664, 16'o000000);
`MEM('o072666, 16'o000000);
`MEM('o072670, 16'o000000);
`MEM('o072672, 16'o000000);
`MEM('o072674, 16'o000000);
`MEM('o072676, 16'o000000);
`MEM('o072700, 16'o000000);
`MEM('o072702, 16'o000000);
`MEM('o072704, 16'o000000);
`MEM('o072706, 16'o000000);
`MEM('o072710, 16'o000000);
`MEM('o072712, 16'o000000);
`MEM('o072714, 16'o000000);
`MEM('o072716, 16'o000000);
`MEM('o072720, 16'o000000);
`MEM('o072722, 16'o000000);
`MEM('o072724, 16'o000000);
`MEM('o072726, 16'o000000);
`MEM('o072730, 16'o000000);
`MEM('o072732, 16'o000000);
`MEM('o072734, 16'o000000);
`MEM('o072736, 16'o000000);
`MEM('o072740, 16'o000000);
`MEM('o072742, 16'o000000);
`MEM('o072744, 16'o000000);
`MEM('o072746, 16'o000000);
`MEM('o072750, 16'o000000);
`MEM('o072752, 16'o000000);
`MEM('o072754, 16'o000000);
`MEM('o072756, 16'o000000);
`MEM('o072760, 16'o000000);
`MEM('o072762, 16'o000000);
`MEM('o072764, 16'o000000);
`MEM('o072766, 16'o000000);
`MEM('o072770, 16'o000000);
`MEM('o072772, 16'o000000);
`MEM('o072774, 16'o000000);
`MEM('o072776, 16'o000000);
`MEM('o073000, 16'o000000);
`MEM('o073002, 16'o000000);
`MEM('o073004, 16'o000000);
`MEM('o073006, 16'o000000);
`MEM('o073010, 16'o000000);
`MEM('o073012, 16'o000000);
`MEM('o073014, 16'o000000);
`MEM('o073016, 16'o000000);
`MEM('o073020, 16'o000000);
`MEM('o073022, 16'o000000);
`MEM('o073024, 16'o000000);
`MEM('o073026, 16'o000000);
`MEM('o073030, 16'o000000);
`MEM('o073032, 16'o000000);
`MEM('o073034, 16'o000000);
`MEM('o073036, 16'o000000);
`MEM('o073040, 16'o000000);
`MEM('o073042, 16'o000000);
`MEM('o073044, 16'o000000);
`MEM('o073046, 16'o000000);
`MEM('o073050, 16'o000000);
`MEM('o073052, 16'o000000);
`MEM('o073054, 16'o000000);
`MEM('o073056, 16'o000000);
`MEM('o073060, 16'o000000);
`MEM('o073062, 16'o000000);
`MEM('o073064, 16'o000000);
`MEM('o073066, 16'o000000);
`MEM('o073070, 16'o000000);
`MEM('o073072, 16'o000000);
`MEM('o073074, 16'o000000);
`MEM('o073076, 16'o000000);
`MEM('o073100, 16'o000000);
`MEM('o073102, 16'o000000);
`MEM('o073104, 16'o000000);
`MEM('o073106, 16'o000000);
`MEM('o073110, 16'o000000);
`MEM('o073112, 16'o000000);
`MEM('o073114, 16'o000000);
`MEM('o073116, 16'o000000);
`MEM('o073120, 16'o000000);
`MEM('o073122, 16'o000000);
`MEM('o073124, 16'o000000);
`MEM('o073126, 16'o000000);
`MEM('o073130, 16'o000000);
`MEM('o073132, 16'o000000);
`MEM('o073134, 16'o000000);
`MEM('o073136, 16'o000000);
`MEM('o073140, 16'o000000);
`MEM('o073142, 16'o000000);
`MEM('o073144, 16'o000000);
`MEM('o073146, 16'o000000);
`MEM('o073150, 16'o000000);
`MEM('o073152, 16'o000000);
`MEM('o073154, 16'o000000);
`MEM('o073156, 16'o000000);
`MEM('o073160, 16'o000000);
`MEM('o073162, 16'o000000);
`MEM('o073164, 16'o000000);
`MEM('o073166, 16'o000000);
`MEM('o073170, 16'o000000);
`MEM('o073172, 16'o000000);
`MEM('o073174, 16'o000000);
`MEM('o073176, 16'o000000);
`MEM('o073200, 16'o000000);
`MEM('o073202, 16'o000000);
`MEM('o073204, 16'o000000);
`MEM('o073206, 16'o000000);
`MEM('o073210, 16'o000000);
`MEM('o073212, 16'o000000);
`MEM('o073214, 16'o000000);
`MEM('o073216, 16'o000000);
`MEM('o073220, 16'o000000);
`MEM('o073222, 16'o000000);
`MEM('o073224, 16'o000000);
`MEM('o073226, 16'o000000);
`MEM('o073230, 16'o000000);
`MEM('o073232, 16'o000000);
`MEM('o073234, 16'o000000);
`MEM('o073236, 16'o000000);
`MEM('o073240, 16'o000000);
`MEM('o073242, 16'o000000);
`MEM('o073244, 16'o000000);
`MEM('o073246, 16'o000000);
`MEM('o073250, 16'o000000);
`MEM('o073252, 16'o000000);
`MEM('o073254, 16'o000000);
`MEM('o073256, 16'o000000);
`MEM('o073260, 16'o000000);
`MEM('o073262, 16'o000000);
`MEM('o073264, 16'o000000);
`MEM('o073266, 16'o000000);
`MEM('o073270, 16'o000000);
`MEM('o073272, 16'o000000);
`MEM('o073274, 16'o000000);
`MEM('o073276, 16'o000000);
`MEM('o073300, 16'o000000);
`MEM('o073302, 16'o000000);
`MEM('o073304, 16'o000000);
`MEM('o073306, 16'o000000);
`MEM('o073310, 16'o000000);
`MEM('o073312, 16'o000000);
`MEM('o073314, 16'o000000);
`MEM('o073316, 16'o000000);
`MEM('o073320, 16'o000000);
`MEM('o073322, 16'o000000);
`MEM('o073324, 16'o000000);
`MEM('o073326, 16'o000000);
`MEM('o073330, 16'o000000);
`MEM('o073332, 16'o000000);
`MEM('o073334, 16'o000000);
`MEM('o073336, 16'o000000);
`MEM('o073340, 16'o000000);
`MEM('o073342, 16'o000000);
`MEM('o073344, 16'o000000);
`MEM('o073346, 16'o000000);
`MEM('o073350, 16'o000000);
`MEM('o073352, 16'o000000);
`MEM('o073354, 16'o000000);
`MEM('o073356, 16'o000000);
`MEM('o073360, 16'o000000);
`MEM('o073362, 16'o000000);
`MEM('o073364, 16'o000000);
`MEM('o073366, 16'o000000);
`MEM('o073370, 16'o000000);
`MEM('o073372, 16'o000000);
`MEM('o073374, 16'o000000);
`MEM('o073376, 16'o000000);
`MEM('o073400, 16'o000000);
`MEM('o073402, 16'o000000);
`MEM('o073404, 16'o000000);
`MEM('o073406, 16'o000000);
`MEM('o073410, 16'o000000);
`MEM('o073412, 16'o000000);
`MEM('o073414, 16'o000000);
`MEM('o073416, 16'o000000);
`MEM('o073420, 16'o000000);
`MEM('o073422, 16'o000000);
`MEM('o073424, 16'o000000);
`MEM('o073426, 16'o000000);
`MEM('o073430, 16'o000000);
`MEM('o073432, 16'o000000);
`MEM('o073434, 16'o000000);
`MEM('o073436, 16'o000000);
`MEM('o073440, 16'o000000);
`MEM('o073442, 16'o000000);
`MEM('o073444, 16'o000000);
`MEM('o073446, 16'o000000);
`MEM('o073450, 16'o000000);
`MEM('o073452, 16'o000000);
`MEM('o073454, 16'o000000);
`MEM('o073456, 16'o000000);
`MEM('o073460, 16'o000000);
`MEM('o073462, 16'o000000);
`MEM('o073464, 16'o000000);
`MEM('o073466, 16'o000000);
`MEM('o073470, 16'o000000);
`MEM('o073472, 16'o000000);
`MEM('o073474, 16'o000000);
`MEM('o073476, 16'o000000);
`MEM('o073500, 16'o000000);
`MEM('o073502, 16'o000000);
`MEM('o073504, 16'o000000);
`MEM('o073506, 16'o000000);
`MEM('o073510, 16'o000000);
`MEM('o073512, 16'o000000);
`MEM('o073514, 16'o000000);
`MEM('o073516, 16'o000000);
`MEM('o073520, 16'o000000);
`MEM('o073522, 16'o000000);
`MEM('o073524, 16'o000000);
`MEM('o073526, 16'o000000);
`MEM('o073530, 16'o000000);
`MEM('o073532, 16'o000000);
`MEM('o073534, 16'o000000);
`MEM('o073536, 16'o000000);
`MEM('o073540, 16'o000000);
`MEM('o073542, 16'o000000);
`MEM('o073544, 16'o000000);
`MEM('o073546, 16'o000000);
`MEM('o073550, 16'o000000);
`MEM('o073552, 16'o000000);
`MEM('o073554, 16'o000000);
`MEM('o073556, 16'o000000);
`MEM('o073560, 16'o000000);
`MEM('o073562, 16'o000000);
`MEM('o073564, 16'o000000);
`MEM('o073566, 16'o000000);
`MEM('o073570, 16'o000000);
`MEM('o073572, 16'o000000);
`MEM('o073574, 16'o000000);
`MEM('o073576, 16'o000000);
`MEM('o073600, 16'o000000);
`MEM('o073602, 16'o000000);
`MEM('o073604, 16'o000000);
`MEM('o073606, 16'o000000);
`MEM('o073610, 16'o000000);
`MEM('o073612, 16'o000000);
`MEM('o073614, 16'o000000);
`MEM('o073616, 16'o000000);
`MEM('o073620, 16'o000000);
`MEM('o073622, 16'o000000);
`MEM('o073624, 16'o000000);
`MEM('o073626, 16'o000000);
`MEM('o073630, 16'o000000);
`MEM('o073632, 16'o000000);
`MEM('o073634, 16'o000000);
`MEM('o073636, 16'o000000);
`MEM('o073640, 16'o000000);
`MEM('o073642, 16'o000000);
`MEM('o073644, 16'o000000);
`MEM('o073646, 16'o000000);
`MEM('o073650, 16'o000000);
`MEM('o073652, 16'o000000);
`MEM('o073654, 16'o000000);
`MEM('o073656, 16'o000000);
`MEM('o073660, 16'o000000);
`MEM('o073662, 16'o000000);
`MEM('o073664, 16'o000000);
`MEM('o073666, 16'o000000);
`MEM('o073670, 16'o000000);
`MEM('o073672, 16'o000000);
`MEM('o073674, 16'o000000);
`MEM('o073676, 16'o000000);
`MEM('o073700, 16'o000000);
`MEM('o073702, 16'o000000);
`MEM('o073704, 16'o000000);
`MEM('o073706, 16'o000000);
`MEM('o073710, 16'o000000);
`MEM('o073712, 16'o000000);
`MEM('o073714, 16'o000000);
`MEM('o073716, 16'o000000);
`MEM('o073720, 16'o000000);
`MEM('o073722, 16'o000000);
`MEM('o073724, 16'o000000);
`MEM('o073726, 16'o000000);
`MEM('o073730, 16'o000000);
`MEM('o073732, 16'o000000);
`MEM('o073734, 16'o000000);
`MEM('o073736, 16'o000000);
`MEM('o073740, 16'o000000);
`MEM('o073742, 16'o000000);
`MEM('o073744, 16'o000000);
`MEM('o073746, 16'o000000);
`MEM('o073750, 16'o000000);
`MEM('o073752, 16'o000000);
`MEM('o073754, 16'o000000);
`MEM('o073756, 16'o000000);
`MEM('o073760, 16'o000000);
`MEM('o073762, 16'o000000);
`MEM('o073764, 16'o000000);
`MEM('o073766, 16'o000000);
`MEM('o073770, 16'o000000);
`MEM('o073772, 16'o000000);
`MEM('o073774, 16'o000000);
`MEM('o073776, 16'o000000);
`MEM('o074000, 16'o000000);
`MEM('o074002, 16'o000000);
`MEM('o074004, 16'o000000);
`MEM('o074006, 16'o000000);
`MEM('o074010, 16'o000000);
`MEM('o074012, 16'o000000);
`MEM('o074014, 16'o000000);
`MEM('o074016, 16'o000000);
`MEM('o074020, 16'o000000);
`MEM('o074022, 16'o000000);
`MEM('o074024, 16'o000000);
`MEM('o074026, 16'o000000);
`MEM('o074030, 16'o000000);
`MEM('o074032, 16'o000000);
`MEM('o074034, 16'o000000);
`MEM('o074036, 16'o000000);
`MEM('o074040, 16'o000000);
`MEM('o074042, 16'o000000);
`MEM('o074044, 16'o000000);
`MEM('o074046, 16'o000000);
`MEM('o074050, 16'o000000);
`MEM('o074052, 16'o000000);
`MEM('o074054, 16'o000000);
`MEM('o074056, 16'o000000);
`MEM('o074060, 16'o000000);
`MEM('o074062, 16'o000000);
`MEM('o074064, 16'o000000);
`MEM('o074066, 16'o000000);
`MEM('o074070, 16'o000000);
`MEM('o074072, 16'o000000);
`MEM('o074074, 16'o000000);
`MEM('o074076, 16'o000000);
`MEM('o074100, 16'o000000);
`MEM('o074102, 16'o000000);
`MEM('o074104, 16'o000000);
`MEM('o074106, 16'o000000);
`MEM('o074110, 16'o000000);
`MEM('o074112, 16'o000000);
`MEM('o074114, 16'o000000);
`MEM('o074116, 16'o000000);
`MEM('o074120, 16'o000000);
`MEM('o074122, 16'o000000);
`MEM('o074124, 16'o000000);
`MEM('o074126, 16'o000000);
`MEM('o074130, 16'o000000);
`MEM('o074132, 16'o000000);
`MEM('o074134, 16'o000000);
`MEM('o074136, 16'o000000);
`MEM('o074140, 16'o000000);
`MEM('o074142, 16'o000000);
`MEM('o074144, 16'o000000);
`MEM('o074146, 16'o000000);
`MEM('o074150, 16'o000000);
`MEM('o074152, 16'o000000);
`MEM('o074154, 16'o000000);
`MEM('o074156, 16'o000000);
`MEM('o074160, 16'o000000);
`MEM('o074162, 16'o000000);
`MEM('o074164, 16'o000000);
`MEM('o074166, 16'o000000);
`MEM('o074170, 16'o000000);
`MEM('o074172, 16'o000000);
`MEM('o074174, 16'o000000);
`MEM('o074176, 16'o000000);
`MEM('o074200, 16'o000000);
`MEM('o074202, 16'o000000);
`MEM('o074204, 16'o000000);
`MEM('o074206, 16'o000000);
`MEM('o074210, 16'o000000);
`MEM('o074212, 16'o000000);
`MEM('o074214, 16'o000000);
`MEM('o074216, 16'o000000);
`MEM('o074220, 16'o000000);
`MEM('o074222, 16'o000000);
`MEM('o074224, 16'o000000);
`MEM('o074226, 16'o000000);
`MEM('o074230, 16'o000000);
`MEM('o074232, 16'o000000);
`MEM('o074234, 16'o000000);
`MEM('o074236, 16'o000000);
`MEM('o074240, 16'o000000);
`MEM('o074242, 16'o000000);
`MEM('o074244, 16'o000000);
`MEM('o074246, 16'o000000);
`MEM('o074250, 16'o000000);
`MEM('o074252, 16'o000000);
`MEM('o074254, 16'o000000);
`MEM('o074256, 16'o000000);
`MEM('o074260, 16'o000000);
`MEM('o074262, 16'o000000);
`MEM('o074264, 16'o000000);
`MEM('o074266, 16'o000000);
`MEM('o074270, 16'o000000);
`MEM('o074272, 16'o000000);
`MEM('o074274, 16'o000000);
`MEM('o074276, 16'o000000);
`MEM('o074300, 16'o000000);
`MEM('o074302, 16'o000000);
`MEM('o074304, 16'o000000);
`MEM('o074306, 16'o000000);
`MEM('o074310, 16'o000000);
`MEM('o074312, 16'o000000);
`MEM('o074314, 16'o000000);
`MEM('o074316, 16'o000000);
`MEM('o074320, 16'o000000);
`MEM('o074322, 16'o000000);
`MEM('o074324, 16'o000000);
`MEM('o074326, 16'o000000);
`MEM('o074330, 16'o000000);
`MEM('o074332, 16'o000000);
`MEM('o074334, 16'o000000);
`MEM('o074336, 16'o000000);
`MEM('o074340, 16'o000000);
`MEM('o074342, 16'o000000);
`MEM('o074344, 16'o000000);
`MEM('o074346, 16'o000000);
`MEM('o074350, 16'o000000);
`MEM('o074352, 16'o000000);
`MEM('o074354, 16'o000000);
`MEM('o074356, 16'o000000);
`MEM('o074360, 16'o000000);
`MEM('o074362, 16'o000000);
`MEM('o074364, 16'o000000);
`MEM('o074366, 16'o000000);
`MEM('o074370, 16'o000000);
`MEM('o074372, 16'o000000);
`MEM('o074374, 16'o000000);
`MEM('o074376, 16'o000000);
`MEM('o074400, 16'o000000);
`MEM('o074402, 16'o000000);
`MEM('o074404, 16'o000000);
`MEM('o074406, 16'o000000);
`MEM('o074410, 16'o000000);
`MEM('o074412, 16'o000000);
`MEM('o074414, 16'o000000);
`MEM('o074416, 16'o000000);
`MEM('o074420, 16'o000000);
`MEM('o074422, 16'o000000);
`MEM('o074424, 16'o000000);
`MEM('o074426, 16'o000000);
`MEM('o074430, 16'o000000);
`MEM('o074432, 16'o000000);
`MEM('o074434, 16'o000000);
`MEM('o074436, 16'o000000);
`MEM('o074440, 16'o000000);
`MEM('o074442, 16'o000000);
`MEM('o074444, 16'o000000);
`MEM('o074446, 16'o000000);
`MEM('o074450, 16'o000000);
`MEM('o074452, 16'o000000);
`MEM('o074454, 16'o000000);
`MEM('o074456, 16'o000000);
`MEM('o074460, 16'o000000);
`MEM('o074462, 16'o000000);
`MEM('o074464, 16'o000000);
`MEM('o074466, 16'o000000);
`MEM('o074470, 16'o000000);
`MEM('o074472, 16'o000000);
`MEM('o074474, 16'o000000);
`MEM('o074476, 16'o000000);
`MEM('o074500, 16'o000000);
`MEM('o074502, 16'o000000);
`MEM('o074504, 16'o000000);
`MEM('o074506, 16'o000000);
`MEM('o074510, 16'o000000);
`MEM('o074512, 16'o000000);
`MEM('o074514, 16'o000000);
`MEM('o074516, 16'o000000);
`MEM('o074520, 16'o000000);
`MEM('o074522, 16'o000000);
`MEM('o074524, 16'o000000);
`MEM('o074526, 16'o000000);
`MEM('o074530, 16'o000000);
`MEM('o074532, 16'o000000);
`MEM('o074534, 16'o000000);
`MEM('o074536, 16'o000000);
`MEM('o074540, 16'o000000);
`MEM('o074542, 16'o000000);
`MEM('o074544, 16'o000000);
`MEM('o074546, 16'o000000);
`MEM('o074550, 16'o000000);
`MEM('o074552, 16'o000000);
`MEM('o074554, 16'o000000);
`MEM('o074556, 16'o000000);
`MEM('o074560, 16'o000000);
`MEM('o074562, 16'o000000);
`MEM('o074564, 16'o000000);
`MEM('o074566, 16'o000000);
`MEM('o074570, 16'o000000);
`MEM('o074572, 16'o000000);
`MEM('o074574, 16'o000000);
`MEM('o074576, 16'o000000);
`MEM('o074600, 16'o000000);
`MEM('o074602, 16'o000000);
`MEM('o074604, 16'o000000);
`MEM('o074606, 16'o000000);
`MEM('o074610, 16'o000000);
`MEM('o074612, 16'o000000);
`MEM('o074614, 16'o000000);
`MEM('o074616, 16'o000000);
`MEM('o074620, 16'o000000);
`MEM('o074622, 16'o000000);
`MEM('o074624, 16'o000000);
`MEM('o074626, 16'o000000);
`MEM('o074630, 16'o000000);
`MEM('o074632, 16'o000000);
`MEM('o074634, 16'o000000);
`MEM('o074636, 16'o000000);
`MEM('o074640, 16'o000000);
`MEM('o074642, 16'o000000);
`MEM('o074644, 16'o000000);
`MEM('o074646, 16'o000000);
`MEM('o074650, 16'o000000);
`MEM('o074652, 16'o000000);
`MEM('o074654, 16'o000000);
`MEM('o074656, 16'o000000);
`MEM('o074660, 16'o000000);
`MEM('o074662, 16'o000000);
`MEM('o074664, 16'o000000);
`MEM('o074666, 16'o000000);
`MEM('o074670, 16'o000000);
`MEM('o074672, 16'o000000);
`MEM('o074674, 16'o000000);
`MEM('o074676, 16'o000000);
`MEM('o074700, 16'o000000);
`MEM('o074702, 16'o000000);
`MEM('o074704, 16'o000000);
`MEM('o074706, 16'o000000);
`MEM('o074710, 16'o000000);
`MEM('o074712, 16'o000000);
`MEM('o074714, 16'o000000);
`MEM('o074716, 16'o000000);
`MEM('o074720, 16'o000000);
`MEM('o074722, 16'o000000);
`MEM('o074724, 16'o000000);
`MEM('o074726, 16'o000000);
`MEM('o074730, 16'o000000);
`MEM('o074732, 16'o000000);
`MEM('o074734, 16'o000000);
`MEM('o074736, 16'o000000);
`MEM('o074740, 16'o000000);
`MEM('o074742, 16'o000000);
`MEM('o074744, 16'o000000);
`MEM('o074746, 16'o000000);
`MEM('o074750, 16'o000000);
`MEM('o074752, 16'o000000);
`MEM('o074754, 16'o000000);
`MEM('o074756, 16'o000000);
`MEM('o074760, 16'o000000);
`MEM('o074762, 16'o000000);
`MEM('o074764, 16'o000000);
`MEM('o074766, 16'o000000);
`MEM('o074770, 16'o000000);
`MEM('o074772, 16'o000000);
`MEM('o074774, 16'o000000);
`MEM('o074776, 16'o000000);
`MEM('o075000, 16'o000000);
`MEM('o075002, 16'o000000);
`MEM('o075004, 16'o000000);
`MEM('o075006, 16'o000000);
`MEM('o075010, 16'o000000);
`MEM('o075012, 16'o000000);
`MEM('o075014, 16'o000000);
`MEM('o075016, 16'o000000);
`MEM('o075020, 16'o000000);
`MEM('o075022, 16'o000000);
`MEM('o075024, 16'o000000);
`MEM('o075026, 16'o000000);
`MEM('o075030, 16'o000000);
`MEM('o075032, 16'o000000);
`MEM('o075034, 16'o000000);
`MEM('o075036, 16'o000000);
`MEM('o075040, 16'o000000);
`MEM('o075042, 16'o000000);
`MEM('o075044, 16'o000000);
`MEM('o075046, 16'o000000);
`MEM('o075050, 16'o000000);
`MEM('o075052, 16'o000000);
`MEM('o075054, 16'o000000);
`MEM('o075056, 16'o000000);
`MEM('o075060, 16'o000000);
`MEM('o075062, 16'o000000);
`MEM('o075064, 16'o000000);
`MEM('o075066, 16'o000000);
`MEM('o075070, 16'o000000);
`MEM('o075072, 16'o000000);
`MEM('o075074, 16'o000000);
`MEM('o075076, 16'o000000);
`MEM('o075100, 16'o000000);
`MEM('o075102, 16'o000000);
`MEM('o075104, 16'o000000);
`MEM('o075106, 16'o000000);
`MEM('o075110, 16'o000000);
`MEM('o075112, 16'o000000);
`MEM('o075114, 16'o000000);
`MEM('o075116, 16'o000000);
`MEM('o075120, 16'o000000);
`MEM('o075122, 16'o000000);
`MEM('o075124, 16'o000000);
`MEM('o075126, 16'o000000);
`MEM('o075130, 16'o000000);
`MEM('o075132, 16'o000000);
`MEM('o075134, 16'o000000);
`MEM('o075136, 16'o000000);
`MEM('o075140, 16'o000000);
`MEM('o075142, 16'o000000);
`MEM('o075144, 16'o000000);
`MEM('o075146, 16'o000000);
`MEM('o075150, 16'o000000);
`MEM('o075152, 16'o000000);
`MEM('o075154, 16'o000000);
`MEM('o075156, 16'o000000);
`MEM('o075160, 16'o000000);
`MEM('o075162, 16'o000000);
`MEM('o075164, 16'o000000);
`MEM('o075166, 16'o000000);
`MEM('o075170, 16'o000000);
`MEM('o075172, 16'o000000);
`MEM('o075174, 16'o000000);
`MEM('o075176, 16'o000000);
`MEM('o075200, 16'o000000);
`MEM('o075202, 16'o000000);
`MEM('o075204, 16'o000000);
`MEM('o075206, 16'o000000);
`MEM('o075210, 16'o000000);
`MEM('o075212, 16'o000000);
`MEM('o075214, 16'o000000);
`MEM('o075216, 16'o000000);
`MEM('o075220, 16'o000000);
`MEM('o075222, 16'o000000);
`MEM('o075224, 16'o000000);
`MEM('o075226, 16'o000000);
`MEM('o075230, 16'o000000);
`MEM('o075232, 16'o000000);
`MEM('o075234, 16'o000000);
`MEM('o075236, 16'o000000);
`MEM('o075240, 16'o000000);
`MEM('o075242, 16'o000000);
`MEM('o075244, 16'o000000);
`MEM('o075246, 16'o000000);
`MEM('o075250, 16'o000000);
`MEM('o075252, 16'o000000);
`MEM('o075254, 16'o000000);
`MEM('o075256, 16'o000000);
`MEM('o075260, 16'o000000);
`MEM('o075262, 16'o000000);
`MEM('o075264, 16'o000000);
`MEM('o075266, 16'o000000);
`MEM('o075270, 16'o000000);
`MEM('o075272, 16'o000000);
`MEM('o075274, 16'o000000);
`MEM('o075276, 16'o000000);
`MEM('o075300, 16'o000000);
`MEM('o075302, 16'o000000);
`MEM('o075304, 16'o000000);
`MEM('o075306, 16'o000000);
`MEM('o075310, 16'o000000);
`MEM('o075312, 16'o000000);
`MEM('o075314, 16'o000000);
`MEM('o075316, 16'o000000);
`MEM('o075320, 16'o000000);
`MEM('o075322, 16'o000000);
`MEM('o075324, 16'o000000);
`MEM('o075326, 16'o000000);
`MEM('o075330, 16'o000000);
`MEM('o075332, 16'o000000);
`MEM('o075334, 16'o000000);
`MEM('o075336, 16'o000000);
`MEM('o075340, 16'o000000);
`MEM('o075342, 16'o000000);
`MEM('o075344, 16'o000000);
`MEM('o075346, 16'o000000);
`MEM('o075350, 16'o000000);
`MEM('o075352, 16'o000000);
`MEM('o075354, 16'o000000);
`MEM('o075356, 16'o000000);
`MEM('o075360, 16'o000000);
`MEM('o075362, 16'o000000);
`MEM('o075364, 16'o000000);
`MEM('o075366, 16'o000000);
`MEM('o075370, 16'o000000);
`MEM('o075372, 16'o000000);
`MEM('o075374, 16'o000000);
`MEM('o075376, 16'o000000);
`MEM('o075400, 16'o000000);
`MEM('o075402, 16'o000000);
`MEM('o075404, 16'o000000);
`MEM('o075406, 16'o000000);
`MEM('o075410, 16'o000000);
`MEM('o075412, 16'o000000);
`MEM('o075414, 16'o000000);
`MEM('o075416, 16'o000000);
`MEM('o075420, 16'o000000);
`MEM('o075422, 16'o000000);
`MEM('o075424, 16'o000000);
`MEM('o075426, 16'o000000);
`MEM('o075430, 16'o000000);
`MEM('o075432, 16'o000000);
`MEM('o075434, 16'o000000);
`MEM('o075436, 16'o000000);
`MEM('o075440, 16'o000000);
`MEM('o075442, 16'o000000);
`MEM('o075444, 16'o000000);
`MEM('o075446, 16'o000000);
`MEM('o075450, 16'o000000);
`MEM('o075452, 16'o000000);
`MEM('o075454, 16'o000000);
`MEM('o075456, 16'o000000);
`MEM('o075460, 16'o000000);
`MEM('o075462, 16'o000000);
`MEM('o075464, 16'o000000);
`MEM('o075466, 16'o000000);
`MEM('o075470, 16'o000000);
`MEM('o075472, 16'o000000);
`MEM('o075474, 16'o000000);
`MEM('o075476, 16'o000000);
`MEM('o075500, 16'o000000);
`MEM('o075502, 16'o000000);
`MEM('o075504, 16'o000000);
`MEM('o075506, 16'o000000);
`MEM('o075510, 16'o000000);
`MEM('o075512, 16'o000000);
`MEM('o075514, 16'o000000);
`MEM('o075516, 16'o000000);
`MEM('o075520, 16'o000000);
`MEM('o075522, 16'o000000);
`MEM('o075524, 16'o000000);
`MEM('o075526, 16'o000000);
`MEM('o075530, 16'o000000);
`MEM('o075532, 16'o000000);
`MEM('o075534, 16'o000000);
`MEM('o075536, 16'o000000);
`MEM('o075540, 16'o000000);
`MEM('o075542, 16'o000000);
`MEM('o075544, 16'o000000);
`MEM('o075546, 16'o000000);
`MEM('o075550, 16'o000000);
`MEM('o075552, 16'o000000);
`MEM('o075554, 16'o000000);
`MEM('o075556, 16'o000000);
`MEM('o075560, 16'o000000);
`MEM('o075562, 16'o000000);
`MEM('o075564, 16'o000000);
`MEM('o075566, 16'o000000);
`MEM('o075570, 16'o000000);
`MEM('o075572, 16'o000000);
`MEM('o075574, 16'o000000);
`MEM('o075576, 16'o000000);
`MEM('o075600, 16'o000000);
`MEM('o075602, 16'o000000);
`MEM('o075604, 16'o000000);
`MEM('o075606, 16'o000000);
`MEM('o075610, 16'o000000);
`MEM('o075612, 16'o000000);
`MEM('o075614, 16'o000000);
`MEM('o075616, 16'o000000);
`MEM('o075620, 16'o000000);
`MEM('o075622, 16'o000000);
`MEM('o075624, 16'o000000);
`MEM('o075626, 16'o000000);
`MEM('o075630, 16'o000000);
`MEM('o075632, 16'o000000);
`MEM('o075634, 16'o000000);
`MEM('o075636, 16'o000000);
`MEM('o075640, 16'o000000);
`MEM('o075642, 16'o000000);
`MEM('o075644, 16'o000000);
`MEM('o075646, 16'o000000);
`MEM('o075650, 16'o000000);
`MEM('o075652, 16'o000000);
`MEM('o075654, 16'o000000);
`MEM('o075656, 16'o000000);
`MEM('o075660, 16'o000000);
`MEM('o075662, 16'o000000);
`MEM('o075664, 16'o000000);
`MEM('o075666, 16'o000000);
`MEM('o075670, 16'o000000);
`MEM('o075672, 16'o000000);
`MEM('o075674, 16'o000000);
`MEM('o075676, 16'o000000);
`MEM('o075700, 16'o000000);
`MEM('o075702, 16'o000000);
`MEM('o075704, 16'o000000);
`MEM('o075706, 16'o000000);
`MEM('o075710, 16'o000000);
`MEM('o075712, 16'o000000);
`MEM('o075714, 16'o000000);
`MEM('o075716, 16'o000000);
`MEM('o075720, 16'o000000);
`MEM('o075722, 16'o000000);
`MEM('o075724, 16'o000000);
`MEM('o075726, 16'o000000);
`MEM('o075730, 16'o000000);
`MEM('o075732, 16'o000000);
`MEM('o075734, 16'o000000);
`MEM('o075736, 16'o000000);
`MEM('o075740, 16'o000000);
`MEM('o075742, 16'o000000);
`MEM('o075744, 16'o000000);
`MEM('o075746, 16'o000000);
`MEM('o075750, 16'o000000);
`MEM('o075752, 16'o000000);
`MEM('o075754, 16'o000000);
`MEM('o075756, 16'o000000);
`MEM('o075760, 16'o000000);
`MEM('o075762, 16'o000000);
`MEM('o075764, 16'o000000);
`MEM('o075766, 16'o000000);
`MEM('o075770, 16'o000000);
`MEM('o075772, 16'o000000);
`MEM('o075774, 16'o000000);
`MEM('o075776, 16'o000000);
`MEM('o076000, 16'o000000);
`MEM('o076002, 16'o000000);
`MEM('o076004, 16'o000000);
`MEM('o076006, 16'o000000);
`MEM('o076010, 16'o000000);
`MEM('o076012, 16'o000000);
`MEM('o076014, 16'o000000);
`MEM('o076016, 16'o000000);
`MEM('o076020, 16'o000000);
`MEM('o076022, 16'o000000);
`MEM('o076024, 16'o000000);
`MEM('o076026, 16'o000000);
`MEM('o076030, 16'o000000);
`MEM('o076032, 16'o000000);
`MEM('o076034, 16'o000000);
`MEM('o076036, 16'o000000);
`MEM('o076040, 16'o000000);
`MEM('o076042, 16'o000000);
`MEM('o076044, 16'o000000);
`MEM('o076046, 16'o000000);
`MEM('o076050, 16'o000000);
`MEM('o076052, 16'o000000);
`MEM('o076054, 16'o000000);
`MEM('o076056, 16'o000000);
`MEM('o076060, 16'o000000);
`MEM('o076062, 16'o000000);
`MEM('o076064, 16'o000000);
`MEM('o076066, 16'o000000);
`MEM('o076070, 16'o000000);
`MEM('o076072, 16'o000000);
`MEM('o076074, 16'o000000);
`MEM('o076076, 16'o000000);
`MEM('o076100, 16'o000000);
`MEM('o076102, 16'o000000);
`MEM('o076104, 16'o000000);
`MEM('o076106, 16'o000000);
`MEM('o076110, 16'o000000);
`MEM('o076112, 16'o000000);
`MEM('o076114, 16'o000000);
`MEM('o076116, 16'o000000);
`MEM('o076120, 16'o000000);
`MEM('o076122, 16'o000000);
`MEM('o076124, 16'o000000);
`MEM('o076126, 16'o000000);
`MEM('o076130, 16'o000000);
`MEM('o076132, 16'o000000);
`MEM('o076134, 16'o000000);
`MEM('o076136, 16'o000000);
`MEM('o076140, 16'o000000);
`MEM('o076142, 16'o000000);
`MEM('o076144, 16'o000000);
`MEM('o076146, 16'o000000);
`MEM('o076150, 16'o000000);
`MEM('o076152, 16'o000000);
`MEM('o076154, 16'o000000);
`MEM('o076156, 16'o000000);
`MEM('o076160, 16'o000000);
`MEM('o076162, 16'o000000);
`MEM('o076164, 16'o000000);
`MEM('o076166, 16'o000000);
`MEM('o076170, 16'o000000);
`MEM('o076172, 16'o000000);
`MEM('o076174, 16'o000000);
`MEM('o076176, 16'o000000);
`MEM('o076200, 16'o000000);
`MEM('o076202, 16'o000000);
`MEM('o076204, 16'o000000);
`MEM('o076206, 16'o000000);
`MEM('o076210, 16'o000000);
`MEM('o076212, 16'o000000);
`MEM('o076214, 16'o000000);
`MEM('o076216, 16'o000000);
`MEM('o076220, 16'o000000);
`MEM('o076222, 16'o000000);
`MEM('o076224, 16'o000000);
`MEM('o076226, 16'o000000);
`MEM('o076230, 16'o000000);
`MEM('o076232, 16'o000000);
`MEM('o076234, 16'o000000);
`MEM('o076236, 16'o000000);
`MEM('o076240, 16'o000000);
`MEM('o076242, 16'o000000);
`MEM('o076244, 16'o000000);
`MEM('o076246, 16'o000000);
`MEM('o076250, 16'o000000);
`MEM('o076252, 16'o000000);
`MEM('o076254, 16'o000000);
`MEM('o076256, 16'o000000);
`MEM('o076260, 16'o000000);
`MEM('o076262, 16'o000000);
`MEM('o076264, 16'o000000);
`MEM('o076266, 16'o000000);
`MEM('o076270, 16'o000000);
`MEM('o076272, 16'o000000);
`MEM('o076274, 16'o000000);
`MEM('o076276, 16'o000000);
`MEM('o076300, 16'o000000);
`MEM('o076302, 16'o000000);
`MEM('o076304, 16'o000000);
`MEM('o076306, 16'o000000);
`MEM('o076310, 16'o000000);
`MEM('o076312, 16'o000000);
`MEM('o076314, 16'o000000);
`MEM('o076316, 16'o000000);
`MEM('o076320, 16'o000000);
`MEM('o076322, 16'o000000);
`MEM('o076324, 16'o000000);
`MEM('o076326, 16'o000000);
`MEM('o076330, 16'o000000);
`MEM('o076332, 16'o000000);
`MEM('o076334, 16'o000000);
`MEM('o076336, 16'o000000);
`MEM('o076340, 16'o000000);
`MEM('o076342, 16'o000000);
`MEM('o076344, 16'o000000);
`MEM('o076346, 16'o000000);
`MEM('o076350, 16'o000000);
`MEM('o076352, 16'o000000);
`MEM('o076354, 16'o000000);
`MEM('o076356, 16'o000000);
`MEM('o076360, 16'o000000);
`MEM('o076362, 16'o000000);
`MEM('o076364, 16'o000000);
`MEM('o076366, 16'o000000);
`MEM('o076370, 16'o000000);
`MEM('o076372, 16'o000000);
`MEM('o076374, 16'o000000);
`MEM('o076376, 16'o000000);
`MEM('o076400, 16'o000000);
`MEM('o076402, 16'o000000);
`MEM('o076404, 16'o000000);
`MEM('o076406, 16'o000000);
`MEM('o076410, 16'o000000);
`MEM('o076412, 16'o000000);
`MEM('o076414, 16'o000000);
`MEM('o076416, 16'o000000);
`MEM('o076420, 16'o000000);
`MEM('o076422, 16'o000000);
`MEM('o076424, 16'o000000);
`MEM('o076426, 16'o000000);
`MEM('o076430, 16'o000000);
`MEM('o076432, 16'o000000);
`MEM('o076434, 16'o000000);
`MEM('o076436, 16'o000000);
`MEM('o076440, 16'o000000);
`MEM('o076442, 16'o000000);
`MEM('o076444, 16'o000000);
`MEM('o076446, 16'o000000);
`MEM('o076450, 16'o000000);
`MEM('o076452, 16'o000000);
`MEM('o076454, 16'o000000);
`MEM('o076456, 16'o000000);
`MEM('o076460, 16'o000000);
`MEM('o076462, 16'o000000);
`MEM('o076464, 16'o000000);
`MEM('o076466, 16'o000000);
`MEM('o076470, 16'o000000);
`MEM('o076472, 16'o000000);
`MEM('o076474, 16'o000000);
`MEM('o076476, 16'o000000);
`MEM('o076500, 16'o000000);
`MEM('o076502, 16'o000000);
`MEM('o076504, 16'o000000);
`MEM('o076506, 16'o000000);
`MEM('o076510, 16'o000000);
`MEM('o076512, 16'o000000);
`MEM('o076514, 16'o000000);
`MEM('o076516, 16'o000000);
`MEM('o076520, 16'o000000);
`MEM('o076522, 16'o000000);
`MEM('o076524, 16'o000000);
`MEM('o076526, 16'o000000);
`MEM('o076530, 16'o000000);
`MEM('o076532, 16'o000000);
`MEM('o076534, 16'o000000);
`MEM('o076536, 16'o000000);
`MEM('o076540, 16'o000000);
`MEM('o076542, 16'o000000);
`MEM('o076544, 16'o000000);
`MEM('o076546, 16'o000000);
`MEM('o076550, 16'o000000);
`MEM('o076552, 16'o000000);
`MEM('o076554, 16'o000000);
`MEM('o076556, 16'o000000);
`MEM('o076560, 16'o000000);
`MEM('o076562, 16'o000000);
`MEM('o076564, 16'o000000);
`MEM('o076566, 16'o000000);
`MEM('o076570, 16'o000000);
`MEM('o076572, 16'o000000);
`MEM('o076574, 16'o000000);
`MEM('o076576, 16'o000000);
`MEM('o076600, 16'o000000);
`MEM('o076602, 16'o000000);
`MEM('o076604, 16'o000000);
`MEM('o076606, 16'o000000);
`MEM('o076610, 16'o000000);
`MEM('o076612, 16'o000000);
`MEM('o076614, 16'o000000);
`MEM('o076616, 16'o000000);
`MEM('o076620, 16'o000000);
`MEM('o076622, 16'o000000);
`MEM('o076624, 16'o000000);
`MEM('o076626, 16'o000000);
`MEM('o076630, 16'o000000);
`MEM('o076632, 16'o000000);
`MEM('o076634, 16'o000000);
`MEM('o076636, 16'o000000);
`MEM('o076640, 16'o000000);
`MEM('o076642, 16'o000000);
`MEM('o076644, 16'o000000);
`MEM('o076646, 16'o000000);
`MEM('o076650, 16'o000000);
`MEM('o076652, 16'o000000);
`MEM('o076654, 16'o000000);
`MEM('o076656, 16'o000000);
`MEM('o076660, 16'o000000);
`MEM('o076662, 16'o000000);
`MEM('o076664, 16'o000000);
`MEM('o076666, 16'o000000);
`MEM('o076670, 16'o000000);
`MEM('o076672, 16'o000000);
`MEM('o076674, 16'o000000);
`MEM('o076676, 16'o000000);
`MEM('o076700, 16'o000000);
`MEM('o076702, 16'o000000);
`MEM('o076704, 16'o000000);
`MEM('o076706, 16'o000000);
`MEM('o076710, 16'o000000);
`MEM('o076712, 16'o000000);
`MEM('o076714, 16'o000000);
`MEM('o076716, 16'o000000);
`MEM('o076720, 16'o000000);
`MEM('o076722, 16'o000000);
`MEM('o076724, 16'o000000);
`MEM('o076726, 16'o000000);
`MEM('o076730, 16'o000000);
`MEM('o076732, 16'o000000);
`MEM('o076734, 16'o000000);
`MEM('o076736, 16'o000000);
`MEM('o076740, 16'o000000);
`MEM('o076742, 16'o000000);
`MEM('o076744, 16'o000000);
`MEM('o076746, 16'o000000);
`MEM('o076750, 16'o000000);
`MEM('o076752, 16'o000000);
`MEM('o076754, 16'o000000);
`MEM('o076756, 16'o000000);
`MEM('o076760, 16'o000000);
`MEM('o076762, 16'o000000);
`MEM('o076764, 16'o000000);
`MEM('o076766, 16'o000000);
`MEM('o076770, 16'o000000);
`MEM('o076772, 16'o000000);
`MEM('o076774, 16'o000000);
`MEM('o076776, 16'o000000);
`MEM('o077000, 16'o000000);
`MEM('o077002, 16'o000000);
`MEM('o077004, 16'o000000);
`MEM('o077006, 16'o000000);
`MEM('o077010, 16'o000000);
`MEM('o077012, 16'o000000);
`MEM('o077014, 16'o000000);
`MEM('o077016, 16'o000000);
`MEM('o077020, 16'o000000);
`MEM('o077022, 16'o000000);
`MEM('o077024, 16'o000000);
`MEM('o077026, 16'o000000);
`MEM('o077030, 16'o000000);
`MEM('o077032, 16'o000000);
`MEM('o077034, 16'o000000);
`MEM('o077036, 16'o000000);
`MEM('o077040, 16'o000000);
`MEM('o077042, 16'o000000);
`MEM('o077044, 16'o000000);
`MEM('o077046, 16'o000000);
`MEM('o077050, 16'o000000);
`MEM('o077052, 16'o000000);
`MEM('o077054, 16'o000000);
`MEM('o077056, 16'o000000);
`MEM('o077060, 16'o000000);
`MEM('o077062, 16'o000000);
`MEM('o077064, 16'o000000);
`MEM('o077066, 16'o000000);
`MEM('o077070, 16'o000000);
`MEM('o077072, 16'o000000);
`MEM('o077074, 16'o000000);
`MEM('o077076, 16'o000000);
`MEM('o077100, 16'o000000);
`MEM('o077102, 16'o000000);
`MEM('o077104, 16'o000000);
`MEM('o077106, 16'o000000);
`MEM('o077110, 16'o000000);
`MEM('o077112, 16'o000000);
`MEM('o077114, 16'o000000);
`MEM('o077116, 16'o000000);
`MEM('o077120, 16'o000000);
`MEM('o077122, 16'o000000);
`MEM('o077124, 16'o000000);
`MEM('o077126, 16'o000000);
`MEM('o077130, 16'o000000);
`MEM('o077132, 16'o000000);
`MEM('o077134, 16'o000000);
`MEM('o077136, 16'o000000);
`MEM('o077140, 16'o000000);
`MEM('o077142, 16'o000000);
`MEM('o077144, 16'o000000);
`MEM('o077146, 16'o000000);
`MEM('o077150, 16'o000000);
`MEM('o077152, 16'o000000);
`MEM('o077154, 16'o000000);
`MEM('o077156, 16'o000000);
`MEM('o077160, 16'o000000);
`MEM('o077162, 16'o000000);
`MEM('o077164, 16'o000000);
`MEM('o077166, 16'o000000);
`MEM('o077170, 16'o000000);
`MEM('o077172, 16'o000000);
`MEM('o077174, 16'o000000);
`MEM('o077176, 16'o000000);
`MEM('o077200, 16'o000000);
`MEM('o077202, 16'o000000);
`MEM('o077204, 16'o000000);
`MEM('o077206, 16'o000000);
`MEM('o077210, 16'o000000);
`MEM('o077212, 16'o000000);
`MEM('o077214, 16'o000000);
`MEM('o077216, 16'o000000);
`MEM('o077220, 16'o000000);
`MEM('o077222, 16'o000000);
`MEM('o077224, 16'o000000);
`MEM('o077226, 16'o000000);
`MEM('o077230, 16'o000000);
`MEM('o077232, 16'o000000);
`MEM('o077234, 16'o000000);
`MEM('o077236, 16'o000000);
`MEM('o077240, 16'o000000);
`MEM('o077242, 16'o000000);
`MEM('o077244, 16'o000000);
`MEM('o077246, 16'o000000);
`MEM('o077250, 16'o000000);
`MEM('o077252, 16'o000000);
`MEM('o077254, 16'o000000);
`MEM('o077256, 16'o000000);
`MEM('o077260, 16'o000000);
`MEM('o077262, 16'o000000);
`MEM('o077264, 16'o000000);
`MEM('o077266, 16'o000000);
`MEM('o077270, 16'o000000);
`MEM('o077272, 16'o000000);
`MEM('o077274, 16'o000000);
`MEM('o077276, 16'o000000);
`MEM('o077300, 16'o000000);
`MEM('o077302, 16'o000000);
`MEM('o077304, 16'o000000);
`MEM('o077306, 16'o000000);
`MEM('o077310, 16'o000000);
`MEM('o077312, 16'o000000);
`MEM('o077314, 16'o000000);
`MEM('o077316, 16'o000000);
`MEM('o077320, 16'o000000);
`MEM('o077322, 16'o000000);
`MEM('o077324, 16'o000000);
`MEM('o077326, 16'o000000);
`MEM('o077330, 16'o000000);
`MEM('o077332, 16'o000000);
`MEM('o077334, 16'o000000);
`MEM('o077336, 16'o000000);
`MEM('o077340, 16'o000000);
`MEM('o077342, 16'o000000);
`MEM('o077344, 16'o000000);
`MEM('o077346, 16'o000000);
`MEM('o077350, 16'o000000);
`MEM('o077352, 16'o000000);
`MEM('o077354, 16'o000000);
`MEM('o077356, 16'o000000);
`MEM('o077360, 16'o000000);
`MEM('o077362, 16'o000000);
`MEM('o077364, 16'o000000);
`MEM('o077366, 16'o000000);
`MEM('o077370, 16'o000000);
`MEM('o077372, 16'o000000);
`MEM('o077374, 16'o000000);
`MEM('o077376, 16'o000000);
`MEM('o077400, 16'o000000);
`MEM('o077402, 16'o000000);
`MEM('o077404, 16'o000000);
`MEM('o077406, 16'o000000);
`MEM('o077410, 16'o000000);
`MEM('o077412, 16'o000000);
`MEM('o077414, 16'o000000);
`MEM('o077416, 16'o000000);
`MEM('o077420, 16'o000000);
`MEM('o077422, 16'o000000);
`MEM('o077424, 16'o000000);
`MEM('o077426, 16'o000000);
`MEM('o077430, 16'o000000);
`MEM('o077432, 16'o000000);
`MEM('o077434, 16'o000000);
`MEM('o077436, 16'o000000);
`MEM('o077440, 16'o000000);
`MEM('o077442, 16'o000000);
`MEM('o077444, 16'o000000);
`MEM('o077446, 16'o000000);
`MEM('o077450, 16'o000000);
`MEM('o077452, 16'o000000);
`MEM('o077454, 16'o000000);
`MEM('o077456, 16'o000000);
`MEM('o077460, 16'o000000);
`MEM('o077462, 16'o000000);
`MEM('o077464, 16'o000000);
`MEM('o077466, 16'o000000);
`MEM('o077470, 16'o000000);
`MEM('o077472, 16'o000000);
`MEM('o077474, 16'o000000);
`MEM('o077476, 16'o000000);
`MEM('o077500, 16'o000000);
`MEM('o077502, 16'o000000);
`MEM('o077504, 16'o000000);
`MEM('o077506, 16'o000000);
`MEM('o077510, 16'o000000);
`MEM('o077512, 16'o000000);
`MEM('o077514, 16'o000000);
`MEM('o077516, 16'o000000);
`MEM('o077520, 16'o000000);
`MEM('o077522, 16'o000000);
`MEM('o077524, 16'o000000);
`MEM('o077526, 16'o000000);
`MEM('o077530, 16'o000000);
`MEM('o077532, 16'o000000);
`MEM('o077534, 16'o000000);
`MEM('o077536, 16'o000000);
`MEM('o077540, 16'o000000);
`MEM('o077542, 16'o000000);
`MEM('o077544, 16'o000000);
`MEM('o077546, 16'o000000);
`MEM('o077550, 16'o000000);
`MEM('o077552, 16'o000000);
`MEM('o077554, 16'o000000);
`MEM('o077556, 16'o000000);
`MEM('o077560, 16'o000000);
`MEM('o077562, 16'o000000);
`MEM('o077564, 16'o000000);
`MEM('o077566, 16'o000000);
`MEM('o077570, 16'o000000);
`MEM('o077572, 16'o000000);
`MEM('o077574, 16'o000000);
`MEM('o077576, 16'o000000);
`MEM('o077600, 16'o000000);
`MEM('o077602, 16'o000000);
`MEM('o077604, 16'o000000);
`MEM('o077606, 16'o000000);
`MEM('o077610, 16'o000000);
`MEM('o077612, 16'o000000);
`MEM('o077614, 16'o000000);
`MEM('o077616, 16'o000000);
`MEM('o077620, 16'o000000);
`MEM('o077622, 16'o000000);
`MEM('o077624, 16'o000000);
`MEM('o077626, 16'o000000);
`MEM('o077630, 16'o000000);
`MEM('o077632, 16'o000000);
`MEM('o077634, 16'o000000);
`MEM('o077636, 16'o000000);
`MEM('o077640, 16'o000000);
`MEM('o077642, 16'o000000);
`MEM('o077644, 16'o000000);
`MEM('o077646, 16'o000000);
`MEM('o077650, 16'o000000);
`MEM('o077652, 16'o000000);
`MEM('o077654, 16'o000000);
`MEM('o077656, 16'o000000);
`MEM('o077660, 16'o000000);
`MEM('o077662, 16'o000000);
`MEM('o077664, 16'o000000);
`MEM('o077666, 16'o000000);
`MEM('o077670, 16'o000000);
`MEM('o077672, 16'o000000);
`MEM('o077674, 16'o000000);
`MEM('o077676, 16'o000000);
`MEM('o077700, 16'o000000);
`MEM('o077702, 16'o000000);
`MEM('o077704, 16'o000000);
`MEM('o077706, 16'o000000);
`MEM('o077710, 16'o000000);
`MEM('o077712, 16'o000000);
`MEM('o077714, 16'o000000);
`MEM('o077716, 16'o000000);
`MEM('o077720, 16'o000000);
`MEM('o077722, 16'o000000);
`MEM('o077724, 16'o000000);
`MEM('o077726, 16'o000000);
`MEM('o077730, 16'o000000);
`MEM('o077732, 16'o000000);
`MEM('o077734, 16'o000000);
`MEM('o077736, 16'o000000);
`MEM('o077740, 16'o000000);
`MEM('o077742, 16'o000000);
`MEM('o077744, 16'o000000);
`MEM('o077746, 16'o000000);
`MEM('o077750, 16'o000000);
`MEM('o077752, 16'o000000);
`MEM('o077754, 16'o000000);
`MEM('o077756, 16'o000000);
`MEM('o077760, 16'o000000);
`MEM('o077762, 16'o000000);
`MEM('o077764, 16'o000000);
`MEM('o077766, 16'o000000);
`MEM('o077770, 16'o000000);
`MEM('o077772, 16'o000000);
`MEM('o077774, 16'o000000);
`MEM('o077776, 16'o000000);
end
