// Bootstrap Loader for Hard Disk
// rom.v
// to be included from the top module at the comple

`define MEM(x, y) {mem_hi[(x)/2], mem_lo[(x)/2]}=y

initial
begin
`MEM('o073700, 16'o012700);
`MEM('o073702, 16'o177472);
`MEM('o073704, 16'o012740);
`MEM('o073706, 16'o000003);
`MEM('o073710, 16'o012740);
`MEM('o073712, 16'o140000);
`MEM('o073714, 16'o012740);
`MEM('o073716, 16'o054000);
`MEM('o073720, 16'o012740);
`MEM('o073722, 16'o176000);
`MEM('o073724, 16'o012740);
`MEM('o073726, 16'o000005);
`MEM('o073730, 16'o105710);
`MEM('o073732, 16'o002376);
`MEM('o073734, 16'o000137);
`MEM('o073736, 16'o054000);
`MEM('o073740, 16'o012700);
`MEM('o073742, 16'o177350);
`MEM('o073744, 16'o005040);
`MEM('o073746, 16'o010040);
`MEM('o073750, 16'o012740);
`MEM('o073752, 16'o000003);
`MEM('o073754, 16'o105710);
`MEM('o073756, 16'o002376);
`MEM('o073760, 16'o005737);
`MEM('o073762, 16'o177350);
`MEM('o073764, 16'o001377);
`MEM('o073766, 16'o112710);
`MEM('o073770, 16'o000005);
`MEM('o073772, 16'o105710);
`MEM('o073774, 16'o002376);
`MEM('o073776, 16'o005007);
`MEM('o074000, 16'o000610);
`MEM('o074002, 16'o003000);
`MEM('o074004, 16'o000400);
`MEM('o074006, 16'o000000);

`MEM('o177570, 16'o173700); // switch register
end
